THERMO
   300.000  600.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2                      N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
CH3               121286C   1H   3          G  0300.00   5000.00  1000.00      1
 2.84405160E+00 6.13797410E-03-2.23034522E-06 3.78516080E-10-2.45215903E-14    2
 1.64378086E+04 5.45269728E+00 2.43044281E+00 1.11240987E-02-1.68022034E-05    3
 1.62182872E-08-5.86495262E-12 1.64237813E+04 6.78979397E+00                   4
C2H6               51090C   2H   6    0    0G   300.000  5000.000 2000.00    0 1
 0.13436084E+02 0.36325546E-02-0.24694586E-06-0.11228470E-09 0.15553612E-13    2
-0.18298318E+05-0.56480824E+02 0.81958778E-01 0.24148658E-01-0.12186742E-04    3
 0.31174958E-08-0.34426783E-12-0.11399086E+05 0.20696499E+02                   4
CH4               121286C   1H   4          G  0300.00   5000.00  1000.00      1
 1.68347883E+00 1.02372356E-02-3.87512864E-06 6.78558487E-10-4.50342312E-14    2
-1.00807871E+04 9.62339497E+00 7.78741479E-01 1.74766835E-02-2.78340904E-05    3
 3.04970804E-08-1.22393068E-11-9.82522852E+03 1.37221947E+01                   4
H                 120186H   1               G  0300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 2.54716270E+04-4.60117638E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 2.54716270E+04-4.60117608E-01                   4
H2                121286H   2               G  0300.00   5000.00  1000.00      1
 2.99142337E+00 7.00064411E-04-5.63382869E-08-9.23157818E-12 1.58275179E-15    2
-8.35033997E+02-1.35511017E+00 3.29812431E+00 8.24944174E-04-8.14301529E-07    3
-9.47543433E-11 4.13487224E-13-1.01252087E+03-3.29409409E+00                   4
CH(S)              71291C   1H   1    0    0G   300.000  3000.000 1000.00    0 1
 0.14872259E+01 0.33000924E-02-0.28411702E-06-0.34383971E-09 0.76660243E-13    2
-0.97217761E+03-0.10147021E+02-0.18660052E+01 0.90233106E-02 0.29339509E-06    3
-0.52555964E-08 0.20409182E-11 0.16202820E+03 0.81504984E+01                   4
C(S,R)             71291C   1    0    0    0G   300.000  3000.000 1000.00    0 1
 0.16900997E+01 0.11069085E-02-0.12616481E-06-0.11996654E-09 0.28811839E-13    2
 0.21028852E+05-0.10340458E+02-0.12628431E+01 0.73135700E-02-0.72650602E-06    3
-0.57274971E-08 0.29829661E-11 0.21889631E+05 0.52818985E+01                   4
CH3(S)             71291C   1H   3    0    0G   300.000  3000.000 1000.00    0 1
 0.22271934E+01 0.64840489E-02-0.50900690E-06-0.66263206E-09 0.14445464E-12    2
 0.72205317E+04-0.13843549E+02-0.23782465E+01 0.14169827E-01 0.60410139E-06    3
-0.75244326E-08 0.28128064E-11 0.87938271E+04 0.11347555E+02                   4
CH2(S)             71291C   1H   2    0    0G   300.000  3000.000 1000.00    0 1
 0.17394471E+01 0.51764320E-02-0.42153641E-06-0.53463645E-09 0.11763388E-12    2
-0.70305313E+04-0.12329198E+02-0.25071146E+01 0.12199585E-01 0.59056043E-06    3
-0.66420434E-08 0.24363521E-11-0.55698042E+04 0.10931940E+02                   4
CH2(S,R)          100191C   1H   2    0    0G   300.000  3000.000 1000.00    0 1
 0.17394471E+01 0.51764320E-02-0.42153641E-06-0.53463645E-09 0.11763388E-12    2
 0.24246523E+05-0.12329198E+02-0.25071146E+01 0.12199585E-01 0.59056043E-06    3
-0.66420434E-08 0.24363521E-11 0.25707254E+05 0.10931940E+02                   4
CH(S,R)            71291C   1H   1    0    0G   300.000  3000.000 1000.00    0 1
 0.14872259E+01 0.33000924E-02-0.28411702E-06-0.34383971E-09 0.76660243E-13    2
 0.15069210E+05-0.10147021E+02-0.18660052E+01 0.90233106E-02 0.29339509E-06    3
-0.52555964E-08 0.20409182E-11 0.16203417E+05 0.81504984E+01                   4
D                  71291C   1    0    0    0G   300.000  3000.000 1000.00    0 1
 0.16900997E+01 0.11069085E-02-0.12616481E-06-0.11996654E-09 0.28811839E-13    2
-0.56464282E+03-0.10340458E+02-0.12628431E+01 0.73135700E-02-0.72650602E-06    3
-0.57274971E-08 0.29829661E-11 0.29613477E+03 0.52818985E+01                   4

END
