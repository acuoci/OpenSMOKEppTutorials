!***********************************************************************
!SURFACE MECHANISM OF THE PARTIAL OXIDATION OF CH4 ON RHODIUM
!***********************************************************************
!****                                                                  *
!****     CPO OF CH4 ON Rh - SURFACE MECHANISM                         *
!****                                                                  *
!****     Version 1.0   February 13, 2001                              *
!****                                                                  *
!****     O. Deutschmann, R. Schwiedernoch, L. Maier,                  *
!****        Heidelberg University, Germany                            *
!****     S. Tummala, L. D. Schmidt, University of Minnesota, USA      *
!****                                                                  *
!****                                                                  *
!****     NOTE: That is a first version that needs further             *
!****           improvements, e.g. methanization, reforming etc.!!!    *
!****                                                                  *
!****                                                                  *
!****     Ref:  O. Deutschmann, R. Schwiedernoch, L.I. Maier,          *
!****           D. Chatterjee. Natural Gas Conversion in Monolithic    *
!****           Catalysts: Interaction of Chemical Reactions and       *
!****           Transport Phenomena.  Natural Gas Conversion VI,       *
!****           Studies in Surface Science and Catalysis 136,          *
!****           E. Iglesia, J.J. Spivey, T.H. Fleisch (eds.),          *
!****           p. 215-258, Elsevier, 2001                             *
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     J/mol  *
!****                                                                  *
!****                                                                  *
!**** SURFACE CHEMKIN format  21.01.06, tested with Vers.4.0.1         *
!****                                                                  *
!***********************************************************************

THERMO
   300.000  1000.000  3000.000
   
H2                121286H   2               G  0300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633828E-06-0.09231578E-10 0.15827519E-14    2
-0.08350340E+04-0.13551101E+01 0.03298124E+02 0.08249441E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.10125209E+04-0.03294094E+02                   4
H                 120186H   1               G  0300.00   5000.00  1000.00      1
 0.02500000E+02 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.02547162E+06-0.04601176E+01 0.02500000E+02 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.02547162E+06-0.04601176E+01                   4
O2                121386O   2               G  0300.00   5000.00  1000.00      1
 0.03697578E+02 0.06135197E-02-0.12588420E-06 0.01775281E-09-0.11364354E-14    2
-0.12339301E+04 0.03189165E+02 0.03212936E+02 0.11274864E-02-0.05756150E-05    3
 0.13138773E-08-0.08768554E-11-0.10052490E+04 0.06034737E+02                   4
O                 120186O   1               G  0300.00   5000.00  1000.00      1
 0.02542059E+02-0.02755061E-03-0.03102803E-07 0.04551067E-10-0.04368051E-14    2
 0.02923080E+06 0.04920308E+02 0.02946428E+02-0.16381665E-02 0.02421031E-04    3
-0.16028431E-08 0.03890696E-11 0.02914764E+06 0.02963995E+02                   4
OH                121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 0.03886888E+05 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 0.03606781E+05 0.13588605E+01                   4
H2O                20387H   2O   1          G  0300.00   5000.00  1000.00      1
 0.02672145E+02 0.03056293E-01-0.08730260E-05 0.12009964E-09-0.06391618E-13    2
-0.02989921E+06 0.06862817E+02 0.03386842E+02 0.03474982E-01-0.06354696E-04    3
 0.06968581E-07-0.02506588E-10-0.03020811E+06 0.02590232E+02                   4
CH4                     C   1H   4          G   300.00   5000.00  1000.00      1
 1.68347883E+00 1.02372356E-02-3.87512864E-06 6.78558487E-10-4.50342312E-14    2
-1.00807871E+04 9.62339497E+00 7.78741479E-01 1.74766835E-02-2.78340904E-05    3
 3.04970804E-08-1.22393068E-11-9.82522852E+03 1.37221947E+01                   4
CO                      C   1O   1          G   300.00   5000.00  1000.00      1
 3.02507806E+00 1.44268852E-03-5.63082779E-07 1.01858133E-10-6.91095156E-15    2
-1.42683496E+04 6.10821772E+00 3.26245165E+00 1.51194085E-03-3.88175522E-06    3
 5.58194424E-09-2.47495123E-12-1.43105391E+04 4.84889698E+00                   4
CO2                     C   1O   2    0     G   300.00   5000.00  1000.00      1
 4.45362282E+00 3.14016873E-03-1.27841054E-06 2.39399667E-10-1.66903319E-14    2
-4.89669609E+04-9.55395877E-01 2.27572465E+00 9.92207229E-03-1.04091132E-05    3
 6.86668678E-09-2.11728009E-12-4.83731406E+04 1.01884880E+01                   4
N2                J 3/77N   20   00   00   0G   300.000  5000.000              1
 0.28532899E+01 0.16022128E-02-0.62936893E-06 0.11441022E-09-0.78057465E-14    2
-0.89008093E+03 0.63964897E+01 0.37044177E+01-0.14218753E-02 0.28670392E-05    3
-0.12028885E-08-0.13954677E-13-0.10640795E+04 0.22336285E+01                   4
AR                L 5/66AR  100  000  000  0G   300.000  5000.000              1
 0.25000000E 01 0.             0.             0.             0.                2
-0.74537502E 03 0.43660006E 01 0.25000000E 01 0.             0.                3
 0.             0.            -0.74537498E 03 0.43660006E 01                   4
 
O(s)               92491O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.19454180E+01 0.91761647E-03-0.11226719E-06-0.99099624E-10 0.24307699E-13    2
-0.14005187E+05-0.11531663E+02-0.94986904E+00 0.74042305E-02-0.10451424E-05    3
-0.61120420E-08 0.33787992E-11-0.13209912E+05 0.36137905E+01                   4
O2(s)              92491O   2Rh  1          I    300.00   3000.00 1000.00      1
 0.35989249E+01 0.20437732E-02-0.23878221E-06-0.22041054E-09 0.53299430E-13    2
-0.41095444E+04-0.21604582E+02-0.20174649E+01 0.14146218E-01-0.16376665E-05    3
-0.11264421E-07 0.60101386E-11-0.25084473E+04 0.79811935E+01                   4
H(s)               92491H   1Rh  1          I    300.00   3000.00 1000.00      1
 0.10696996E+01 0.15432230E-02-0.15500922E-06-0.16573165E-09 0.38359347E-13    2
-0.50546128E+04-0.71555238E+01-0.13029877E+01 0.54173199E-02 0.31277972E-06    3
-0.32328533E-08 0.11362820E-11-0.42277075E+04 0.58743238E+01                   4
H2(s)              92491H   2Rh  1          I    300.00   3000.00 1000.00      1
 0.15330955E+01 0.34586885E-02-0.32622225E-06-0.36824219E-09 0.83855205E-13    2
-0.36401533E+04-0.10822206E+02-0.21517782E+01 0.87039210E-02 0.11154106E-05    3
-0.42477102E-08 0.96133203E-12-0.22640681E+04 0.97397461E+01                   4
H2O(s)             92491O   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.25803051E+01 0.49570827E-02-0.46894056E-06-0.52633137E-09 0.11998322E-12    2
-0.38302234E+05-0.17406322E+02-0.27651553E+01 0.13315115E-01 0.10127695E-05    3
-0.71820083E-08 0.22813776E-11-0.36398055E+05 0.12098145E+02                   4
OH(s)              92491O   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.18249973E+01 0.32501565E-02-0.31197541E-06-0.34603206E-09 0.79171472E-13    2
-0.26685492E+05-0.12280891E+02-0.20340881E+01 0.93662683E-02 0.66275214E-06    3
-0.52074887E-08 0.17088735E-11-0.25319949E+05 0.89863186E+01                   4
Rh(s)                   Rh  1               S    300.0    3000.0  1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(s)                  0C   1O   1Rh  1     S    300.00   3000.00 1000.00      1
 0.47083778E+01 0.96037297E-03-0.11805279E-06-0.76883826E-10 0.18232000E-13    2
-0.32311723E+05-0.16719593E+02 0.48907466E+01 0.68134235E-04 0.19768814E-06    3
 0.12388669E-08-0.90339249E-12-0.32297836E+05-0.17453161E+02                   4
CO2(s)            081292C   1O   2Rh  1     I   300.00   3000.00  1000.00      1
 0.46900000E+00 0.62660000E-02 0.00000000E-00 0.00000000E-00 0.00000000E-00    2
-0.50458700E+05-0.45550000E+01 0.46900000E+00 0.62662000E-02 0.00000000E-00    3
 0.00000000E-00 0.00000000E-00-0.50458700E+05-0.45550000E+01                   4
C(s)                   0C   1Rh  1          I    300.00   3000.00 1000.00      1
 0.15792824E+01 0.36528701E-03-0.50657672E-07-0.34884855E-10 0.88089699E-14    2
 0.99535752E+04-0.30240495E+01 0.58924019E+00 0.25012842E-02-0.34229498E-06    3
-0.18994346E-08 0.10190406E-11 0.10236923E+05 0.21937017E+01                   4
CH(s)                  0C   1H   1Rh  1     I    300.00   3000.00 1000.00      1
-0.48242472E-02 0.30446239E-02-0.16066099E-06-0.29041700E-09 0.57999924E-13    2
 0.22595219E+05 0.56677818E+01 0.84157485E+00 0.13095380E-02 0.28464575E-06    3
 0.63862904E-09-0.42766658E-12 0.22332801E+05 0.11452305E+01                   4
CH2(s)                 0C   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.74076122E+00 0.48032533E-02-0.32825633E-06-0.47779786E-09 0.10073452E-12    2
 0.10443752E+05 0.40842086E+00-0.14876404E+00 0.51396289E-02 0.11211075E-05    3
-0.82755452E-09-0.44572345E-12 0.10878700E+05 0.57451882E+01                   4
CH3(s)                 0C   1H   3Rh  1     I    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
HCO(s)                 0C   1H   1O   1Rh  1S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
CH4(s)                 0C   1H   4Rh  1     I    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4

O_Rh                    O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
O2(s)                   O   2Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H_Rh                    H   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2(s)                   H   2Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O_Rh                  O   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
OH_Rh                   O   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
_Rh_                    Rh  1               S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO_Rh                   C   1O   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO2_Rh                  C   1O   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C_Rh                    C   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH_Rh                   C   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH2_Rh                  C   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH3_Rh                  C   1H   3Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH4_Rh                  C   1H   4Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
