THERMO
  300.0   1000.0   3000.0
Rh(s)                   Rh  1               S    300.0    3000.0  1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
O(s)               92491O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H(s)               92491H   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
OH(s)              92491O   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O(s)             92491O   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(s)                  0C   1O   1Rh  1     S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO2(s)            081292C   1O   2Rh  1     S   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C(s)                   0C   1Rh  1          S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH(s)                  0C   1H   1Rh  1     S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH2(s)                 0C   1H   2Rh  1     S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH3(s)                 0C   1H   3Rh  1     S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
COOH(s)                0C   1H   1O   2Rh  1S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
HCOO(s)                0C   1H   1O   2Rh  2S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2                      H   2               G    300.00   5000.00 1000.00      1
 .299142220E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033546E+03-.135510641E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
O2                      O   2               G    300.00   5000.00 1000.00      1
 .369757685E+01 .613519690E-03-.125884200E-06 .177528100E-10-.113643500E-14    2
-.123392966E+04 .318917125E+01 .321293600E+01 .112748610E-02-.575614990E-06    3
 .131387700E-08-.876855390E-12-.100524900E+04 .603473900E+01                   4
H2O               L 8/89H   2O   1          G 200.000  3500.000  1000.000      1
 3.03399249E+00 2.17691804E-03-1.64072518E-07-9.70419870E-11 1.68200992E-14    2
-3.00042971E+04 4.96677010E+00 4.19864056E+00-2.03643410E-03 6.52040211E-06    3
-5.48797062E-09 1.77197817E-12-3.02937267E+04-8.49032208E-01                   4
H                 L 7/88H   1               G 200.000  3500.000  1000.000      1
 2.50000001E+00-2.30842973E-11 1.61561948E-14-4.73515235E-18 4.98197357E-22    2
 2.54736599E+04-4.46682914E-01 2.50000000E+00 7.05332819E-13-1.99591964E-15    3
 2.30081632E-18-9.27732332E-22 2.54736599E+04-4.46682853E-01                   4
OH                RUS 78O   1H   1          G 200.000  3500.000  1000.000      1
 3.09288767E+00 5.48429716E-04 1.26505228E-07-8.79461556E-11 1.17412376E-14    2
 3.85865700E+03 4.47669610E+00 3.99201543E+00-2.40131752E-03 4.61793841E-06    3
-3.88113333E-09 1.36411470E-12 3.61508056E+03-1.03925458E-01                   4
O                       O   1               G    300.00   5000.00 1000.00      1
 2.56942078E+00-8.59741137E-05 4.19484589E-08-1.00177799E-11 1.22833691E-15    2
 2.92175791E+04 4.78433864E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3
-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00                   4
HCOO              T04/97H   1C   1O   2     G 298.150  5000.000  1000.000      1
 5.97791811E+00 3.24247847E-03-1.46666291E-06 2.91808902E-10-2.10704956E-14    2
-2.04910217E+04-7.12854015E+00-3.01936623E+01 2.54607495E-01-6.43484728E-04    3
 6.92943698E-07-2.65871657E-10-1.59887826E+04 1.47958586E+02-1.81158000E+04    4
COOH              RUS 79H   1C   1O   2     G 200.000  6000.000  1000.000      1
 0.53920264E+01 0.41122622E-02-0.14819726E-05 0.23988016E-09-0.14390635E-13    2
-0.27670863E+05-0.22350810E+01 0.29220825E+01 0.76245184E-02 0.32988630E-05    3
-0.10713524E-07 0.51158655E-11-0.26838359E+05 0.11292583E+02-0.25617866E+05    4
CO                TPIS79C   1O   1          G 200.000  3500.000  1000.000      1
 2.71518561E+00 2.06252743E-03-9.98825771E-07 2.30053008E-10-2.03647716E-14    2
-1.41518724E+04 7.81868772E+00 3.57953347E+00-6.10353680E-04 1.01681433E-06    3
 9.07005884E-10-9.04424499E-13-1.43440860E+04 3.50840928E+00                   4
CO2               L 7/88C   1O   2          G 200.000  3500.000  1000.000      1
 3.85746029E+00 4.41437026E-03-2.21481404E-06 5.23490188E-10-4.72084164E-14    2
-4.87591660E+04 2.27163806E+00 2.35677352E+00 8.98459677E-03-7.12356269E-06    3
 2.45919022E-09-1.43699548E-13-4.83719697E+04 9.90105222E+00                   4
C                 L11/88C   1               G 200.000  3500.000  1000.000      1
 2.49266888E+00 4.79889284E-05-7.24335020E-08 3.74291029E-11-4.87277893E-15    2
 8.54512953E+04 4.80150373E+00 2.55423955E+00-3.21537724E-04 7.33792245E-07    3
-7.32234889E-10 2.66521446E-13 8.54438832E+04 4.53130848E+00                   4
CH                TPIS79C   1H   1          G 200.000  3500.000  1000.000      1
 2.87846473E+00 9.70913681E-04 1.44445655E-07-1.30687849E-10 1.76079383E-14    2
 7.10124364E+04 5.48497999E+00 3.48981665E+00 3.23835541E-04-1.68899065E-06    3
 3.16217327E-09-1.40609067E-12 7.07972934E+04 2.08401108E+00                   4
CH2               L S/93C   1H   2          G 200.000  3500.000  1000.000      1
 2.87410113E+00 3.65639292E-03-1.40894597E-06 2.60179549E-10-1.87727567E-14    2
 4.62636040E+04 6.17119324E+00 3.76267867E+00 9.68872143E-04 2.79489841E-06    3
-3.85091153E-09 1.68741719E-12 4.60040401E+04 1.56253185E+00                   4
CH3               L11/89C   1H   3          G 200.000  3500.000  1000.000      1
 2.28571772E+00 7.23990037E-03-2.98714348E-06 5.95684644E-10-4.67154394E-14    2
 1.67755843E+04 8.48007179E+00 3.67359040E+00 2.01095175E-03 5.73021856E-06    3
-6.87117425E-09 2.54385734E-12 1.64449988E+04 1.60456433E+00                   4
CH4               L 8/88C   1H   4          G 200.000  3500.000  1000.000      1
 7.48514950E-02 1.33909467E-02-5.73285809E-06 1.22292535E-09-1.01815230E-13    2
-9.46834459E+03 1.84373180E+01 5.14987613E+00-1.36709788E-02 4.91800599E-05    3
-4.84743026E-08 1.66693956E-11-1.02466476E+04-4.64130376E+00                   4
N2                      N   2               G    300.00   5000.00 1000.00      1
 .292663788E+01 .148797700E-02-.568476030E-06 .100970400E-09-.675335090E-14    2
-.922795384E+03 .598054018E+01 .329867700E+01 .140823990E-02-.396322180E-05    3
 .564151480E-08-.244485400E-11-.102090000E+04 .395037200E+01                   4
C3H8              120186C   3H   8          G   300.000  5000.000 1000.00      1
 7.52521700e+00 1.88903400e-02-6.28392400e-06 9.17937300e-10-4.81241000e-14    2
-1.64645500e+04-1.78439000e+01 8.96920800e-01 2.66898600e-02 5.43142500e-06    3
-2.12600100e-08 9.24333000e-12-1.39549200e+04 1.93553300e+01                   4
C3H6              120186C   3H   6          G   300.000  5000.000 1000.00      1
 6.73225700e+00 1.49083400e-02-4.94989900e-06 7.21202200e-10-3.76620400e-14    2
-9.23570300e+02-1.33133500e+01 1.49330700e+00 2.09251800e-02 4.48679400e-06    3
-1.66891200e-08 7.15814600e-12 1.07482600e+03 1.61453400e+01                   4
HE                      HE  1               G    300.00   5000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
-.745375000E+03 .928723974E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375000E+03 .928723974E+00                   4
AR                      AR  1               G    300.00   5000.00 1000.00      1
 .312500009E+01-.140625050E-02 .937500490E-06-.156250080E-09 .000000000E+00    2
-.940687583E+03 .103823694E+01 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375100E+03 .436600100E+01                   4
N2                      N   2               G    300.00   5000.00 1000.00      1
 .292663788E+01 .148797700E-02-.568476030E-06 .100970400E-09-.675335090E-14    2
-.922795384E+03 .598054018E+01 .329867700E+01 .140823990E-02-.396322180E-05    3
 .564151480E-08-.244485400E-11-.102090000E+04 .395037200E+01                   4
NO                      O   1N   1          G    300.00   5000.00 1000.00      1
 .324543589E+01 .126913800E-02-.501589000E-06 .916928270E-10-.627541890E-14    2
 .980084032E+04 .641728767E+01 .337654100E+01 .125306300E-02-.330275000E-05    3
 .521781020E-08-.244626190E-11 .981796100E+04 .582959200E+01                   4
N2O                     O   1N   2          G    300.00   5000.00 1000.00      1
 .471897567E+01 .287371290E-02-.119749600E-05 .225055100E-09-.157533690E-13    2
 .816581343E+04-.165723704E+01 .254305700E+01 .949219330E-02-.979277500E-05    3
 .626384410E-08-.190182510E-11 .876510200E+04 .951122400E+01                   4
O2                      O   2               G    300.00   5000.00 1000.00      1
 .369757685E+01 .613519690E-03-.125884200E-06 .177528100E-10-.113643500E-14    2
-.123392966E+04 .318917125E+01 .321293600E+01 .112748610E-02-.575614990E-06    3
 .131387700E-08-.876855390E-12-.100524900E+04 .603473900E+01                   4
NO2                     O   2N   1          G    300.00   5000.00 1000.00      1
 .468285677E+01 .246242900E-02-.104225900E-05 .197690200E-09-.139171700E-13    2
 .226129300E+04 .988610659E+00 .267060000E+01 .783849970E-02-.806386380E-05    3
 .616171380E-08-.232014990E-11 .289629000E+04 .116120700E+02                   4
HNO                     H   1O   1N   1     G    300.00   5000.00 1000.00      1
 .361514436E+01 .321248500E-02-.126033690E-05 .226729700E-09-.153623600E-13    2
 .106619122E+05 .481025325E+01 .278440200E+01 .660964610E-02-.930022270E-05    3
 .943798020E-08-.375314580E-11 .109187800E+05 .903562900E+01                   4
HNNO                    H   1O   1N   2     G    300.00   5000.00 1500.00      1
 .699121930E+01 .187597000E-02-.212458400E-06-.671047200E-10 .123050800E-13    2
 .249756641E+05-.112352384E+02 .223829800E+01 .135920000E-01-.117987300E-04    3
 .539297100E-08-.101085900E-11 .266025900E+05 .141367900E+02                   4
HNO2                    H   1O   2N   1     G    300.00   5000.00 1500.00      1
 .647962840E+01 .199527400E-02-.174038700E-06-.969587200E-10 .170148000E-13    2
-.999926943E+04-.106728455E+02 .193483800E+01 .101003600E-01-.496461600E-05    3
 .870112000E-09-.232413500E-14-.810548400E+04 .147325000E+02                   4
HONO                    H   1O   2N   1     G    300.00   5000.00 1000.00      1
 .548688978E+01 .421806500E-02-.164914300E-05 .297187700E-09-.202114800E-13    2
-.112686489E+05-.299698546E+01 .229041300E+01 .140992200E-01-.136787200E-04    3
 .749878000E-08-.187690500E-11-.104319500E+05 .132807700E+02                   4
HONO2                   H   1O   3N   1     G    300.00   5000.00 1500.00      1
 .975613289E+01 .190094800E-02-.324002000E-06-.397663900E-10 .110033400E-13    2
-.194224157E+05-.269001236E+02 .787766800E+00 .238232900E-01-.220596400E-04    3
 .103404800E-07-.197285700E-11-.163044200E+05 .210896400E+02                   4
H2                      H   2               G    300.00   5000.00 1000.00      1
 .299142220E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033546E+03-.135510641E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
N2H2                    H   2N   2          G    300.00   5000.00 1000.00      1
 .337118994E+01 .603996800E-02-.230385300E-05 .406278900E-09-.271314400E-13    2
 .241817095E+05 .498055769E+01 .161799940E+01 .130631220E-01-.171571100E-04    3
 .160560790E-07-.609363800E-11 .246752600E+05 .137946700E+02                   4
H2O                     H   2O   1          G    300.00   5000.00 1000.00      1
 .267214569E+01 .305629290E-02-.873026070E-06 .120099600E-09-.639161790E-14    2
-.298992115E+05 .686281125E+01 .338684200E+01 .347498200E-02-.635469590E-05    3
 .696858040E-08-.250658800E-11-.302081100E+05 .259023200E+01                   4
H2O2                    H   2O   2          G    300.00   5000.00 1000.00      1
 .457316594E+01 .433613590E-02-.147468900E-05 .234890300E-09-.143165410E-13    2
-.180069531E+05 .501137915E+00 .338875300E+01 .656922580E-02-.148501200E-06    3
-.462580510E-08 .247151410E-11-.176631400E+05 .678536300E+01                   4
NH3                     H   3N   1          G    300.00   5000.00 1000.00      1
 .246189456E+01 .605916650E-02-.200497610E-05 .313600310E-09-.193831700E-13    2
-.649326483E+04 .747215046E+01 .220435100E+01 .101147600E-01-.146526500E-04    3
 .144723500E-07-.532850890E-11-.652548900E+04 .812714000E+01                   4
N2H4                    H   4N   2          G    300.00   5000.00 1000.00      1
 .497732211E+01 .959551900E-02-.354763900E-05 .612429900E-09-.402979500E-13    2
 .934121983E+04-.296302077E+01 .644260600E-01 .274973000E-01-.289945100E-04    3
 .174524000E-07-.442228200E-11 .104519200E+05 .212778900E+02                   4
CO                      C   1O   1          G    300.00   5000.00 1000.00      1
 .302507617E+01 .144268900E-02-.563082720E-06 .101858100E-09-.691095110E-14    2
-.142683499E+05 .610822521E+01 .326245100E+01 .151194100E-02-.388175520E-05    3
 .558194380E-08-.247495100E-11-.143105400E+05 .484889700E+01                   4
CO2                     C   1O   2          G    300.00   5000.00 1000.00      1
 .445362582E+01 .314016800E-02-.127841100E-05 .239399610E-09-.166903300E-13    2
-.489669524E+05-.955420007E+00 .227572400E+01 .992207230E-02-.104091100E-04    3
 .686668590E-08-.211728010E-11-.483731400E+05 .101884900E+02                   4
HCN                     C   1H   1N   1     G    300.00   5000.00 1000.00      1
 .365007798E+01 .346099790E-02-.127427900E-05 .221765490E-09-.147717700E-13    2
 .149839102E+05 .239321426E+01 .249046200E+01 .861127950E-02-.103103400E-04    3
 .748149810E-08-.222910900E-11 .152083400E+05 .790498000E+01                   4
HNCO                    C   1H   1O   1N   1G    300.00   5000.00 1000.00      1
 .621186395E+01 .229713690E-02-.221612790E-06-.122204400E-09 .227240590E-13    2
-.147707257E+05-.801661658E+01 .369405900E+01 .665723530E-02-.505446810E-07    3
-.347341090E-08 .136056900E-11-.139197600E+05 .571273900E+01                   4
HCNO                    C   1H   1O   1N   1G    300.00   5000.00 1000.00      1
 .669241213E+01 .236836030E-02-.237151000E-06-.127550300E-09 .240713700E-13    2
 .169473623E+05-.124543537E+02 .318485800E+01 .975231640E-02-.128020300E-05    3
-.616310380E-08 .322627490E-11 .179790700E+05 .612384200E+01                   4
HOCN                    C   1H   1O   1N   1G    300.00   5000.00 1000.00      1
 .564560836E+01 .229820610E-02-.216262900E-06-.121480100E-09 .223863610E-13    2
-.317811025E+04-.359027798E+01 .362829200E+01 .566418420E-02-.117020600E-06    3
-.234863800E-08 .801640220E-12-.247592500E+04 .747682300E+01                   4
CH2O                    C   1H   2O   1     G    300.00   5000.00 1000.00      1
 .299560858E+01 .668132120E-02-.262895400E-05 .473715290E-09-.321251710E-13    2
-.153203666E+05 .691256052E+01 .165273100E+01 .126314400E-01-.188816790E-04    3
 .205003110E-07-.841323710E-11-.148654000E+05 .137848200E+02                   4
HCO3H                   C   1H   2O   3     G    300.00   5000.00 1378.00      1
 .987503581E+01 .464663708E-02-.167230522E-05 .268624413E-09-.159595232E-13    2
-.380502456E+05-.224938942E+02 .242464726E+01 .219706380E-01-.168705546E-04    3
 .625612194E-08-.911645843E-12-.354828006E+05 .175027796E+02                   4
CH3NO                   C   1H   3O   1N   1G    300.00   5000.00 1500.00      1
 .882055478E+01 .370623300E-02-.289474100E-06-.189791000E-09 .323754400E-13    2
 .536285603E+04-.221322539E+02 .210995500E+01 .151782200E-01-.707178900E-05    3
 .151061100E-08-.160420400E-12 .829361200E+04 .156970200E+02                   4
CH3NO2                  C   1H   3O   2N   1G    300.00   5000.00 1382.00      1
 .750407068E+01 .952121946E-02-.327760562E-05 .508678596E-09-.294455378E-13    2
-.121591399E+05-.115088778E+02-.370775080E+00 .283702793E-01-.208339624E-04    3
 .808980673E-08-.130521082E-11-.945681543E+04 .306459151E+02                   4
CH3ONO                  C   1H   3O   2N   1G    300.00   5000.00 1500.00      1
 .113612738E+02 .415934900E-02-.414567000E-06-.169514000E-09 .302873200E-13    2
-.128147952E+05-.354542296E+02 .149034500E+01 .264543300E-01-.211233200E-04    3
 .941439900E-08-.181120500E-11-.912578200E+04 .181376600E+02                   4
CH3ONO2                 C   1H   3O   3N   1G    300.00   5000.00 1500.00      1
 .143618741E+02 .411224300E-02-.511305200E-06-.149643600E-09 .301215600E-13    2
-.197243835E+05-.513183467E+02 .780335400E+00 .345420400E-01-.282232800E-04    3
 .123232400E-07-.230216400E-11-.146534600E+05 .224575200E+02                   4
CH4                     C   1H   4          G    300.00   5000.00 1000.00      1
 .168346564E+01 .102372400E-01-.387512820E-05 .678558490E-09-.450342310E-13    2
-.100807773E+05 .962347575E+01 .778741700E+00 .174766800E-01-.278340900E-04    3
 .304970800E-07-.122393100E-10-.982522800E+04 .137221900E+02                   4
CH3OH                   C   1H   4O   1     G    300.00   5000.00 1000.00      1
 .402907793E+01 .937659290E-02-.305025380E-05 .435879300E-09-.222472310E-13    2
-.261579223E+05 .237808255E+01 .266011500E+01 .734150780E-02 .717005010E-05    3
-.879319370E-08 .239056990E-11-.253534800E+05 .112326300E+02                   4
CH3OOH                  C   1H   4O   2     G    300.00   5000.00 1000.00      1
 .563694993E+01 .111814780E-01-.369593390E-05 .407189810E-09 .000000000E+00    2
-.180442749E+05-.124166637E+01 .586865100E+01 .107942400E-01-.364552990E-05    3
 .541291180E-09-.289684390E-13-.181268900E+05-.251762300E+01                   4
C2H2                    C   2H   2          G    300.00   5000.00 1000.00      1
 .443677300E+01 .537603910E-02-.191281610E-05 .328637890E-09-.215670900E-13    2
 .256676622E+05-.280035722E+01 .201356200E+01 .151904500E-01-.161631910E-04    3
 .907899180E-08-.191274600E-11 .261244400E+05 .880537800E+01                   4
CH2CO                   C   2H   2O   1     G    300.00   5000.00 1000.00      1
 .603885318E+01 .580484000E-02-.192095400E-05 .279448500E-09-.145886800E-13    2
-.858343402E+04-.765782305E+01 .297497100E+01 .121187100E-01-.234504600E-05    3
-.646668500E-08 .390564900E-11-.763263700E+04 .867355300E+01                   4
CH3CN                   C   2H   3N   1     G    300.00   5000.00 1000.00      1
 .239240386E+01 .156188730E-01-.791204970E-05 .193723330E-08-.186119560E-12    2
 .849993803E+04 .111452402E+02 .251975310E+01 .135675230E-01-.257640770E-05    3
-.308939670E-08 .142886920E-11 .855337620E+04 .109208680E+02                   4
C2H4                    C   2H   4          G    300.00   5000.00 1000.00      1
 .352841648E+01 .114851800E-01-.441838480E-05 .784460000E-09-.526684780E-13    2
 .442829030E+04 .223039249E+01-.861487900E+00 .279616190E-01-.338867690E-04    3
 .278515200E-07-.973787890E-11 .557304700E+04 .242114800E+02                   4
C2H4O                   C   2H   4O   1     G    300.00   5000.00 1000.00      1
 .385543260E+01 .146081760E-01-.526121540E-05 .628115500E-09 .000000000E+00    2
-.851874300E+04 .214156911E+01-.130385500E+01 .282461720E-01-.170593430E-04    3
 .394753470E-08 .000000000E+00-.707559900E+04 .289352600E+02                   4
CH3CHO                  C   2H   4O   1     G    300.00   5000.00 1000.00      1
 .586869116E+01 .107942400E-01-.364552990E-05 .541291180E-09-.289684390E-13    2
-.226457128E+05-.601321650E+01 .250569500E+01 .133699100E-01 .467195290E-05    3
-.112814000E-07 .426356610E-11-.212458800E+05 .133508900E+02                   4
CH3COOH                 C   2H   4O   2     G    300.00   5000.00 1000.00      1
 .691666936E+01 .128920800E-01-.420990320E-05 .458049540E-09 .000000000E+00    2
-.553508487E+05-.102392103E+02 .846928500E+00 .292145000E-01-.186455200E-04    3
 .464098720E-08 .000000000E+00-.536761800E+05 .211901500E+02                   4
CH3OCHO                 C   2H   4O   2     G    300.00   5000.00 1686.00      1
 .869123518E+01 .115503122E-01-.427782486E-05 .702533059E-09-.424333552E-13    2
-.464364769E+05-.189301478E+02 .308839783E+01 .203760048E-01-.684777040E-05    3
-.728186203E-09 .562130216E-12-.441855167E+05 .125364719E+02                   4
C2-OQOOH                C   2H   4O   3     G    300.00   5000.00 1380.00      1
 .124064339E+02 .947233784E-02-.328107928E-05 .513772211E-09-.299872803E-13    2
-.349123142E+05-.339479874E+02 .552382546E+01 .242068306E-01-.152898974E-04    3
 .501728362E-08-.696406358E-12-.323406789E+05 .357240645E+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   5000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
DME-OQOOH               C   2H   4O   4     G    300.00   5000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
C2H6                    C   2H   6          G    300.00   5000.00 1000.00      1
 .482597579E+01 .138404300E-01-.455725790E-05 .672496720E-09-.359816110E-13    2
-.127178296E+05-.523976258E+01 .146253900E+01 .154946700E-01 .578050690E-05    3
-.125783200E-07 .458626710E-11-.112391800E+05 .144322900E+02                   4
C2H5OH                  C   2H   6O   1     G    300.00   5000.00 1000.00      1
 .434717120E+01 .186288000E-01-.677946700E-05 .816592600E-09 .000000000E+00    2
-.306615743E+05 .324247304E+01 .576535800E+00 .289451200E-01-.161002000E-04    3
 .359164100E-08 .000000000E+00-.296359500E+05 .227081300E+02                   4
CH3OCH3                 C   2H   6O   1     G    300.00   5000.00 1368.00      1
 .827732656E+01 .132135539E-01-.453264362E-05 .705316507E-09-.409933283E-13    2
-.261980897E+05-.215181376E+02 .150763450E+01 .239914228E-01-.868910500E-05    3
-.966835762E-10 .489319361E-12-.232810894E+05 .167317297E+02                   4
C2H5OOH                 C   2H   6O   2     G    300.00   5000.00 1000.00      1
 .914611907E+01 .144611400E-01-.455120020E-05 .475780030E-09 .000000000E+00    2
-.236690607E+05-.205899250E+02 .223998300E+01 .310914290E-01-.170933710E-04    3
 .329379790E-08 .000000000E+00-.216018500E+05 .158174300E+02                   4
C3H2                    C   3H   2          G    300.00   5000.00 1000.00      1
 .767099642E+01 .274874900E-02-.437094300E-06-.645559900E-10 .166388700E-13    2
 .625972092E+05-.123689926E+02 .316671400E+01 .248257200E-01-.459163700E-04    3
 .426801900E-07-.148215200E-10 .635042100E+05 .886944600E+01                   4
PC3H4                   C   3H   4          G    300.00   5000.00 1000.00      1
 .281460543E+01 .185524496E-01-.955026768E-05 .239951370E-08-.237485257E-12    2
 .207010771E+05 .860604972E+01 .146175323E+01 .246026602E-01-.190219395E-04    3
 .860363422E-08-.166729240E-11 .209209793E+05 .149262585E+02                   4
AC3H4                   C   3H   4          G    300.00   5000.00 1400.07      1
 .977625145E+01 .530213820E-02-.370111790E-06-.302638610E-09 .508958110E-13    2
 .195497314E+05-.307705909E+02 .253983090E+01 .163343700E-01-.176495000E-05    3
-.464736520E-08 .172913110E-11 .225124300E+05 .993570230E+01                   4
C2H3CHO                 C   3H   4O   1     G    300.00   5000.00 1393.00      1
 .104184607E+02 .948963321E-02-.329310529E-05 .516279203E-09-.301587291E-13    2
-.149629790E+05-.307232511E+02 .292355162E+00 .354321417E-01-.294936324E-04    3
 .128100124E-07-.226144108E-11-.116521584E+05 .228878280E+02                   4
C3H6                    C   3H   6          G    300.00   5000.00 1000.00      1
 .673231663E+01 .149083400E-01-.494989900E-05 .721202210E-09-.376620390E-13    2
-.923623057E+03-.133137684E+02 .149330700E+01 .209251700E-01 .448679380E-05    3
-.166891190E-07 .715814600E-11 .107482600E+04 .161453400E+02                   4
C2H5CHO                 C   3H   6O   1     G    300.00   5000.00 1378.00      1
 .102429148E+02 .139641989E-01-.476248001E-05 .738105706E-09-.427759503E-13    2
-.274145137E+05-.285357348E+02 .216308444E+01 .295501264E-01-.152446252E-04    3
 .349503947E-08-.238896627E-12-.242260137E+05 .161153348E+02                   4
C3H5OH                  C   3H   6O   1     G    300.00   5000.00 1000.00      1
 .665875100E+01 .179008100E-01-.612801520E-05 .983706560E-09-.609475850E-13    2
-.187194550E+05-.446185680E+01 .332545570E+01 .251539630E-01-.163055650E-04    3
 .121609030E-07-.500807290E-11-.174250940E+05 .139104030E+02                   4
CH3COCH3                C   3H   6O   1     G    300.00   5000.00 1374.00      1
 .991426580E+01 .146030709E-01-.506085765E-05 .792682855E-09-.462739645E-13    2
-.311168055E+05-.286116537E+02 .130767163E+01 .292021742E-01-.119045617E-04    3
 .652150087E-09 .467751203E-12-.275328269E+05 .196395025E+02                   4
C3H6O                   C   3H   6O   1     G    300.00   5000.00 1000.00      1
 .433142310E+01 .236433890E-01-.875060690E-05 .106889830E-08 .000000000E+00    2
-.138496111E+05 .215169726E+01 .507423500E+00 .318789710E-01-.137497700E-04    3
 .165647900E-08 .000000000E+00-.126239100E+05 .226350900E+02                   4
C3H5OOH                 C   3H   6O   2     G    300.00   5000.00 1382.00      1
 .139268456E+02 .135384067E-01-.474335693E-05 .748389157E-09-.439105886E-13    2
-.132537727E+05-.456757848E+02 .221491505E+01 .390935107E-01-.258809564E-04    3
 .870894601E-08-.120793929E-11-.896037969E+04 .179425329E+02                   4
C3-OQOOH                C   3H   6O   3     G    300.00   5000.00 1391.00      1
 .170285271E+02 .130716784E-01-.459310856E-05 .726135156E-09-.426658337E-13    2
-.416334217E+05-.592513577E+02 .768933034E+00 .546905880E-01-.465072405E-04    3
 .203159585E-07-.358398999E-11-.363238861E+05 .268291637E+02                   4
C3H8                    C   3H   8          G    300.00   5000.00 1000.00      1
 .752530602E+01 .188903400E-01-.628392400E-05 .917937280E-09-.481240960E-13    2
-.164646226E+05-.178445202E+02 .896921000E+00 .266898590E-01 .543142510E-05    3
-.212600000E-07 .924333010E-11-.139549200E+05 .193553300E+02                   4
IC3H7OH                 C   3H   8O   1     G    300.00   5000.00 1000.00      1
 .577239007E+01 .268947430E-01-.111795290E-04 .211392460E-08-.149320990E-12    2
-.361710675E+05-.384089810E+01-.176838920E+00 .452559560E-01-.319190720E-04    3
 .123062880E-07-.201412540E-11-.346643940E+05 .263322250E+02                   4
NC3H7OH                 C   3H   8O   1     G    300.00   5000.00 1396.00      1
 .107520626E+02 .180260472E-01-.603049401E-05 .922166246E-09-.529319319E-13    2
-.361555719E+05-.310977038E+02 .978207214E-01 .420500918E-01-.267066894E-04    3
 .903941170E-08-.128324751E-11-.323437836E+05 .264700804E+02                   4
C3H7OOH                 C   3H   8O   2     G    300.00   5000.00 1388.00      1
 .150655849E+02 .170865595E-01-.593183927E-05 .930136673E-09-.543384935E-13    2
-.301371140E+05-.515057998E+02 .783525746E+00 .504826223E-01-.365089942E-04    3
 .140377750E-07-.226737156E-11-.251105573E+05 .253041175E+02                   4
C4H2                    C   4H   2          G    300.00   5000.00 1000.00      1
 .903147468E+01 .604725210E-02-.194878790E-05 .275486300E-09-.138560800E-13    2
 .529472934E+05-.238511290E+02 .400519100E+01 .198100000E-01-.986587660E-05    3
-.663515820E-08 .607741290E-11 .542406400E+05 .184573600E+01                   4
C4H4                    C   4H   4          G    300.00   5000.00 1000.00      1
 .665080310E+01 .161294300E-01-.719388700E-05 .149817800E-08-.118641100E-12    2
 .311958636E+05-.979559836E+01-.191524700E+01 .527508700E-01-.716559400E-04    3
 .550724200E-07-.172862200E-10 .329785000E+05 .314199800E+02                   4
C4H6                    C   4H   6          G    300.00   5000.00 1000.00      1
 .823794980E+01 .173695890E-01-.615923200E-05 .979908060E-09-.578075590E-13    2
 .923259930E+04-.203418190E+02 .112443850E+00 .343711770E-01-.111106630E-04    3
-.921096660E-08 .620841700E-11 .118022620E+05 .230917180E+02                   4
IC3H5CHO                C   4H   6O   1     G    300.00   5000.00 1396.00      1
 .136175682E+02 .137917192E-01-.473370118E-05 .736655226E-09-.420097974E-13    2
-.199994281E+05-.472987367E+02 .627183793E+00 .466780254E-01-.374430631E-04    3
 .158330542E-07-.273952155E-11-.157203117E+05 .216034294E+02                   4
MACRIL                  C   4H   6O   2     G    300.00   5000.00 1000.00      1
 .962595080E+01 .202069860E-01-.684948550E-05 .109063620E-08-.671284990E-13    2
-.414857110E+05-.177414250E+02-.929250120E+00 .565245670E-01-.531143270E-04    3
 .263405850E-07-.484636380E-11-.390243280E+05 .347643170E+02                   4
IC4H8                   C   4H   8          G    300.00   5000.00 1388.00      1
 .112258330E+02 .181795798E-01-.620348592E-05 .961444458E-09-.557088057E-13    2
-.769983777E+04-.373306704E+02 .938433173E+00 .390547287E-01-.216437148E-04    3
 .587267077E-08-.614435479E-12-.374817891E+04 .191442985E+02                   4
NC4H8                   C   4H   8          G    300.00   5000.00 1000.00      1
 .205358410E+01 .343505070E-01-.158831970E-04 .330896620E-08-.253610450E-12    2
-.213972310E+04 .155432010E+02 .118113800E+01 .308533800E-01 .508652470E-05    3
-.246548880E-07 .111101930E-10-.179040040E+04 .210624690E+02                   4
C3H7CHO                 C   4H   8O   1     G    300.00   5000.00 1000.00      1
 .885754490E+01 .242627260E-01-.846559850E-05 .137561310E-08-.858588980E-13    2
-.294816840E+05-.174775160E+02 .666312930E+00 .477311800E-01-.329931100E-04    3
 .121733550E-07-.165405020E-11-.272346390E+05 .246936170E+02                   4
MEK                     C   4H   8O   1     G    300.00   5000.00 1000.00      1
 .929655016E+01 .229172746E-01-.822048591E-05 .132404838E-08-.791751980E-13    2
-.334442311E+05-.204993263E+02 .661978185E+01 .851847835E-02 .510322077E-04    3
-.658433042E-07 .249110484E-10-.315251691E+05-.109485469E+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   5000.00 1391.00      1
 .137503148E+02 .183126722E-01-.628572629E-05 .978250756E-09-.568538653E-13    2
-.326938845E+05-.477281342E+02-.273021382E+00 .489696307E-01-.312770049E-04    3
 .100052945E-07-.127512074E-11-.276054737E+05 .283451139E+02                   4
C4H7OH                  C   4H   8O   1     G    300.00   5000.00 1000.00      1
 .863167950E+01 .241150480E-01-.832957180E-05 .134433130E-08-.835340300E-13    2
-.230779140E+05-.163015210E+02 .173864090E+01 .369849060E-01-.680297030E-05    3
-.128647340E-07 .662652570E-11-.209184180E+05 .207395880E+02                   4
C4H8O                   C   4H   8O   1     G    300.00   5000.00 1371.00      1
 .154228514E+02 .170211052E-01-.606347951E-05 .967354762E-09-.571992419E-13    2
-.220196123E+05-.613882135E+02-.253690104E+01 .543995707E-01-.343390305E-04    3
 .101079922E-07-.110262736E-11-.152980680E+05 .367400719E+02                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   5000.00 1390.00      1
 .195047991E+02 .181701803E-01-.634838146E-05 .999797067E-09-.585883751E-13    2
-.450007951E+05-.705122130E+02 .549934041E+00 .642751153E-01-.501779820E-04    3
 .203546231E-07-.338767418E-11-.385647626E+05 .307013051E+02                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   5000.00 1388.00      1
 .195955254E+02 .180568312E-01-.629994700E-05 .991157547E-09-.580382406E-13    2
-.461054913E+05-.709333761E+02 .243440296E+01 .605409309E-01-.481250984E-04    3
 .203656751E-07-.357059537E-11-.402872220E+05 .205488821E+02                   4
NC4H10                  C   4H  10          G    300.00   5000.00 1000.00      1
 .105251152E+02 .235908740E-01-.785389060E-05 .114561140E-08-.599309560E-13    2
-.204952316E+05-.321928008E+02 .157641510E+01 .345897230E-01 .697016090E-05    3
-.281636370E-07 .123751170E-10-.171470040E+05 .178727420E+02                   4
IC4H10                  C   4H  10          G    300.00   5000.00 1000.00      1
 .508434390E+01 .331851280E-01-.124047670E-04 .152753620E-08 .000000000E+00    2
-.195243797E+05-.392308050E+01-.128398800E+01 .519486400E-01-.308267920E-04    3
 .755438110E-08 .000000000E+00-.179038400E+05 .285063500E+02                   4
TC4H9OH                 C   4H  10O   1     G    300.00   5000.00 1395.00      1
 .151183592E+02 .214941230E-01-.730928419E-05 .113021881E-08-.653833962E-13    2
-.450124898E+05-.575375902E+02-.861795957E+00 .603867730E-01-.445191256E-04    3
 .177406426E-07-.295852901E-11-.395611057E+05 .278278048E+02                   4
N1C4H9OH                C   4H  10O   1     G    300.00   5000.00 1389.00      1
 .146461472E+02 .217370421E-01-.745243572E-05 .115877769E-08-.672987557E-13    2
-.406432319E+05-.509926617E+02 .129085275E+00 .529074664E-01-.325907761E-04    3
 .102723019E-07-.133027252E-11-.352672374E+05 .280463660E+02                   4
IC4H9OH                 C   4H  10O   1     G    300.00   5000.00 1426.00      1
 .145203606E+02 .218826590E-01-.741886985E-05 .114493281E-08-.661481541E-13    2
-.415815847E+05-.516504190E+02-.808654483E+00 .568695746E-01-.379891888E-04    3
 .133635469E-07-.195588405E-11-.361485459E+05 .310126347E+02                   4
N2C4H9OH                C   4H  10O   1     G    300.00   5000.00 1390.00      1
 .151582366E+02 .215048627E-01-.741631184E-05 .115764678E-08-.674130532E-13    2
-.429113728E+05-.549620416E+02-.304705097E+00 .567446943E-01-.387293873E-04    3
 .141775813E-07-.220696859E-11-.373601662E+05 .285520284E+02                   4
C4H9OOH                 C   4H  10O   2     G    300.00   5000.00 1389.00      1
 .182257559E+02 .215996217E-01-.748424942E-05 .117205153E-08-.684096331E-13    2
-.342341151E+05-.670536388E+02 .607792497E+00 .624669916E-01-.444490375E-04    3
 .167754668E-07-.265938189E-11-.280070327E+05 .278025473E+02                   4
CYC5H4O                 C   5H   4O   1     G    300.00   5000.00 1000.00      1
 .558734350E+01 .254149730E-01-.929145880E-05 .112347330E-08 .000000000E+00    2
 .339172461E+04-.552979995E+01-.427809100E+01 .546170700E-01-.380993520E-04    3
 .105947040E-07 .000000000E+00 .589093400E+04 .446629800E+02                   4
CYC5H6                  C   5H   6          G    300.00   5000.00 1000.00      1
 .230537462E+00 .409571826E-01-.241588958E-04 .679763480E-08-.736374421E-12    2
 .143779465E+05 .202551234E+02-.513691194E+01 .606953453E-01-.460552837E-04    3
 .128457201E-07 .741214852E-12 .153675713E+05 .461567559E+02                   4
CYC5H8                  C   5H   8          G    300.00   5000.00 1000.00      1
 .772447728E+01 .283223160E-01-.115452360E-04 .215408150E-08-.150541780E-12    2
-.782614232E+03-.197696844E+02 .268981400E+01 .209545500E-02 .113036870E-03    3
-.154080700E-06 .627636580E-10 .231396630E+04 .152940560E+02                   4
C5H8                    C   5H   8          G    300.00   5000.00 1000.00      1
 .797205310E+01 .268614160E-01-.956546320E-05 .113079120E-08 .000000000E+00    2
 .510466811E+04-.185090870E+02 .176636500E+01 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .684030700E+04 .137180600E+02                   4
C5H8O                   C   5H   8O   1     G    300.00   5000.00 1000.00      1
 .154011002E+02 .203490440E-01-.699742510E-05 .109031908E-08-.634192782E-13    2
-.910076428E+04-.580710041E+02-.514624016E+01 .722177875E-01-.580157542E-04    3
 .242093068E-07-.410120178E-11-.236133441E+04 .508920452E+02                   4
MCROT                   C   5H   8O   2     G    300.00   5000.00 1000.00      1
 .110840220E+02 .266681570E-01-.910298150E-05 .145819250E-08-.902072000E-13    2
-.461868520E+05-.238654710E+02 .115411390E+01 .550597160E-01-.356332020E-04    3
 .867407750E-08 .746845670E-12-.435806950E+05 .269868980E+02                   4
C5EN-OQOOH-53           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-54           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-45           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
ETMB583                 C   5H   8O   3     G    300.00   5000.00 1000.00      1
 .164044820E+02 .257082970E-01-.901921340E-05 .147114070E-08-.920586850E-13    2
-.622657890E+05-.550660710E+02-.249091940E+01 .790685040E-01-.564648800E-04    3
 .115540360E-07 .278656790E-11-.573317190E+05 .417407460E+02                   4
C5EN-OQOOH-34           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-43           C   5H   8O   3     G    300.00   5000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
KEHYMB                  C   5H   8O   5     G    300.00   5000.00 1000.00      1
 .130410150E+02 .302430520E-01-.103682550E-04 .166520830E-08-.103159200E-12    2
-.605793360E+05-.352927630E+02-.187604440E+01 .779613480E-01-.656695630E-04    3
 .280818550E-07-.405575270E-11-.569013010E+05 .398655930E+02                   4
NC5H10                  C   5H  10          G    300.00   5000.00 1389.00      1
 .141108203E+02 .228348272E-01-.778626835E-05 .120627491E-08-.698795983E-13    2
-.114335029E+05-.501593461E+02-.541560551E+00 .539629918E-01-.323508738E-04    3
 .977416037E-08-.118534668E-11-.598606169E+04 .297142748E+02                   4
IC5H10                  C   5H  10          G    300.00   5000.00 1000.00      1
 .124808598E+02 .240088830E-01-.777773490E-05 .119128510E-08-.709457860E-13    2
-.864177347E+04-.392940217E+02-.599261880E+00 .540460090E-01-.294562720E-04    3
 .525642110E-08 .585451010E-12-.450159910E+04 .303432560E+02                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   5000.00 1406.00      1
 .182053093E+02 .222888126E-01-.759419141E-05 .117633164E-08-.681511068E-13    2
-.260973639E+05-.785614741E+02-.704702259E+01 .864172552E-01-.702610933E-04    3
 .290540959E-07-.480586102E-11-.179483330E+05 .550571499E+02                   4
NC5H10-O                C   5H  10O   1     G    300.00   5000.00 1373.00      1
 .187152768E+02 .216122625E-01-.768638433E-05 .122492227E-08-.723734176E-13    2
-.274341627E+05-.786690289E+02-.351633623E+01 .686975884E-01-.446579237E-04    3
 .140670556E-07-.174934766E-11-.191663581E+05 .425589840E+02                   4
C4H9CHO                 C   5H  10O   1     G    300.00   5000.00 1381.00      1
 .167965264E+02 .225684519E-01-.767631588E-05 .118769369E-08-.687545554E-13    2
-.356826220E+05-.609064044E+02 .159663472E+01 .543541416E-01-.321020651E-04    3
 .935773559E-08-.106688932E-11-.299841025E+05 .221281498E+02                   4
MB                      C   5H  10O   2     G    300.00   5000.00 1380.00      1
 .190094725E+02 .236503722E-01-.822978452E-05 .129246265E-08-.755862836E-13    2
-.634989152E+05-.732469099E+02 .316208825E+01 .552915358E-01-.311610102E-04    3
 .842394129E-08-.872222021E-12-.573385240E+05 .139723817E+02                   4
MTBE-O                  C   5H  10O   2     G    300.00   5000.00 1397.00      1
 .193844587E+02 .224929046E-01-.748169734E-05 .114123661E-08-.654437288E-13    2
-.558416627E+05-.795832532E+02-.518049059E+01 .839546669E-01-.663790553E-04    3
 .267623941E-07-.432034827E-11-.478415885E+05 .506953652E+02                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   5000.00 1397.00      1
 .237028187E+02 .215843890E-01-.747470111E-05 .117038715E-08-.683143724E-13    2
-.509464263E+05-.948314143E+02 .101097520E+01 .753376897E-01-.559848192E-04    3
 .210040666E-07-.316727025E-11-.432003697E+05 .266737910E+02                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   5000.00 1389.00      1
 .227422860E+02 .225948063E-01-.786379640E-05 .123514506E-08-.722413862E-13    2
-.501979972E+05-.864068664E+02 .227305950E+01 .724929431E-01-.560597536E-04    3
 .231254746E-07-.397203084E-11-.431866364E+05 .229745558E+02                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   5000.00 1386.00      1
 .259492704E+02 .217762181E-01-.754080079E-05 .118109778E-08-.689663912E-13    2
-.659884236E+05-.102260628E+03 .215705064E+01 .770950997E-01-.562944956E-04    3
 .205751475E-07-.301215733E-11-.577585957E+05 .255153989E+02                   4
NC5H12                  C   5H  12          G    300.00   5000.00 1000.00      1
 .142233709E+02 .264253600E-01-.834599270E-05 .125651470E-08-.740004510E-13    2
-.247106388E+05-.503994927E+02-.393634560E+00 .578781330E-01-.285392090E-04    3
 .347472500E-08 .106523800E-11-.198713480E+05 .281908260E+02                   4
NEOC5H12                C   5H  12          G    300.00   5000.00 1397.00      1
 .174488013E+02 .245462377E-01-.835182479E-05 .129219708E-08-.747942850E-13    2
-.292378530E+05-.754164601E+02-.288372771E+01 .722417687E-01-.511106166E-04    3
 .187342407E-07-.280628313E-11-.222171069E+05 .336765462E+02                   4
MTBE                    C   5H  12O   1     G    300.00   5000.00 1000.00      1
 .888656643E+01 .420057870E-01-.178904220E-04 .345077750E-08-.247674430E-12    2
-.405353691E+05-.208281992E+02-.162610860E+01 .742240170E-01-.539682020E-04    3
 .210023490E-07-.342702090E-11-.378579060E+05 .325557600E+02                   4
NC5H11OOH               C   5H  12O   2     G    300.00   5000.00 1391.00      1
 .215962451E+02 .259122865E-01-.896302814E-05 .140202940E-08-.817685827E-13    2
-.395542326E+05-.852046644E+02-.443227141E+00 .781363104E-01-.573273118E-04    3
 .222802059E-07-.361215684E-11-.318952281E+05 .330316890E+02                   4
C6H2                    C   6H   2          G    300.00   5000.00 1000.00      1
 .127565190E+02 .803438100E-02-.261821500E-05 .372506000E-09-.187885000E-13    2
 .807546900E+05-.404126200E+02 .575108500E+01 .263671900E-01-.116675960E-04    3
-.107144980E-07 .879029700E-11 .826201200E+05-.433553200E+01                   4
C6H4                    C   6H   4          G    300.00   5000.00 1000.00      1
 .171831170E+02 .664876580E-02-.124162630E-05 .146974480E-09-.913980130E-14    2
 .550769540E+05-.644351830E+02 .193231390E+01 .390321830E-01-.692271090E-05    3
-.270933570E-07 .157302520E-10 .596919480E+05 .165160230E+02                   4
BENZYNE                 C   6H   4          G    300.00   5000.00 1000.00      1
 .105707063E+02 .156860613E-01-.568267148E-05 .922956737E-09-.554966417E-13    2
 .504976657E+05-.332563927E+02 .721604591E+00 .247976151E-01 .316372209E-04    3
-.653230986E-07 .296082142E-10 .539797980E+05 .216733825E+02                   4
C6H4O2                  C   6H   4O   2     G    300.00   5000.00 1000.00      1
 .148186534E+02 .176963450E-01-.512229240E-05 .482867020E-09 .000000000E+00    2
-.210645982E+05-.499092297E+02-.357739600E+01 .669980650E-01-.485375860E-04    3
 .129924900E-07 .000000000E+00-.159750500E+05 .454022300E+02                   4
LC6H6                   C   6H   6          G    300.00   5000.00 1000.00      1
 .133755312E+02 .181053970E-01-.671790940E-05 .114930710E-08-.753903640E-13    2
 .353349989E+05-.436278915E+02-.284372350E+01 .754240600E-01-.877316710E-04    3
 .551440390E-07-.141557690E-10 .392169020E+05 .371208190E+02                   4
C6H6                    C   6H   6          G    300.00   5000.00 1000.00      1
 .129109067E+02 .172329600E-01-.502421020E-05 .589349680E-09-.194752100E-13    2
 .366437279E+04-.500281184E+02-.313801200E+01 .472310300E-01-.296220700E-05    3
-.326281900E-07 .171869100E-10 .889003000E+04 .365757300E+02                   4
C6H5OH                  C   6H   6O   1     G    300.00   5000.00 1000.00      1
 .141552427E+02 .199350340E-01-.718219540E-05 .116229002E-08-.697147483E-13    2
-.181287441E+05-.517984911E+02-.290978575E+00 .408562397E-01 .242829425E-04    3
-.714477617E-07 .346002146E-10-.134129780E+05 .268745637E+02                   4
MCPTD                   C   6H   8          G    300.00   5000.00 1399.00      1
 .154352848E+02 .199801707E-01-.680270423E-05 .105349633E-08-.610336727E-13    2
 .447456576E+04-.636393642E+02-.665320026E+01 .744640477E-01-.582864186E-04    3
 .231603543E-07-.369017129E-11 .117669311E+05 .538162769E+02                   4
CYC6H8                  C   6H   8          G    300.00   5000.00 1384.00      1
 .167797183E+02 .200748305E-01-.710732570E-05 .112925397E-08-.665827513E-13    2
 .222453062E+04-.729120687E+02-.719572313E+01 .780676798E-01-.620002183E-04    3
 .253310854E-07-.423684696E-11 .104082650E+05 .552451233E+02                   4
CYC6H10                 C   6H  10          G    300.00   5000.00 1388.00      1
 .164687940E+02 .250464584E-01-.873323457E-05 .137353265E-08-.804138942E-13    2
-.977694533E+04-.696690108E+02-.607599781E+01 .751138370E-01-.506516889E-04    3
 .171683701E-07-.235089637E-11-.166592755E+04 .523699408E+02                   4
C6H10-ONE               C   6H  10O   1     G    300.00   5000.00 1382.00      1
 .189587175E+02 .263606964E-01-.929344737E-05 .147257311E-08-.866645349E-13    2
-.391424596E+05-.835594309E+02-.541298687E+01 .749581025E-01-.429010347E-04    3
 .103686234E-07-.655858987E-12-.298390440E+05 .503037294E+02                   4
C5H9CHO                 C   6H  10O   1     G    300.00   5000.00 1369.00      1
 .194648486E+02 .257619052E-01-.914519168E-05 .145563936E-08-.859339746E-13    2
-.393988116E+05-.858349504E+02-.528503736E+01 .742084262E-01-.414393902E-04    3
 .926068588E-08-.391839791E-12-.298547201E+05 .504370563E+02                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   5000.00 1381.00      1
 .208569012E+02 .251723586E-01-.898344923E-05 .143508332E-08-.849382249E-13    2
-.384586302E+05-.102070819E+03-.138345764E+02 .100994913E+00-.688346635E-04    3
 .212451763E-07-.229797219E-11-.260978348E+05 .857505804E+02                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   5000.00 1384.00      1
 .209040427E+02 .249694592E-01-.887525958E-05 .141404459E-08-.835397954E-13    2
-.281106427E+05-.100684615E+03-.120242065E+02 .974927920E-01-.669797836E-04    3
 .211938876E-07-.242310206E-11-.164176421E+05 .774198780E+02                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   5000.00 1388.00      1
 .211309516E+02 .245922161E-01-.870218393E-05 .138238722E-08-.815033630E-13    2
-.270082298E+05-.100017882E+03-.102441734E+02 .947119743E-01-.662992744E-04    3
 .218368996E-07-.269065692E-11-.159562249E+05 .693449458E+02                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   5000.00 1416.00      1
 .160913887E+02 .291196520E-01-.940602358E-05 .140488615E-08-.793370497E-13    2
-.378857796E+05-.754185099E+02-.107476916E+02 .986835275E-01-.783513685E-04    3
 .322824282E-07-.532533650E-11-.294335398E+05 .659825481E+02                   4
ALDEST                  C   6H  10O   3     G    300.00   5000.00 1384.00      1
 .212949599E+02 .266487791E-01-.898035403E-05 .137511216E-08-.789865729E-13    2
-.762788357E+05-.785214726E+02 .521237801E+01 .613142880E-01-.373337900E-04    3
 .119679719E-07-.162337383E-11-.703135588E+05 .903341827E+01                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   5000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   5000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.696293762E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .532148412E+02                   4
CYC6H12                 C   6H  12          G    300.00   5000.00 1373.00      1
 .190852614E+02 .283866516E-01-.999547753E-05 .158256182E-08-.930877430E-13    2
-.260770569E+05-.880292959E+02-.782903355E+01 .809375102E-01-.439655186E-04    3
 .871887784E-08-.486950162E-15-.157787533E+05 .600472718E+02                   4
NC6H12                  C   6H  12          G    300.00   5000.00 1000.00      1
 .186637886E+02 .209714510E-01-.310828090E-05-.686516180E-09 .160236080E-12    2
-.135910200E+05-.708905467E+02 .196862030E+01 .476562310E-01 .660153730E-05    3
-.371481730E-07 .169224630E-10-.771187890E+04 .208592300E+02                   4
ETBE                    C   6H  14O   1     G    300.00   5000.00 1000.00      1
 .107600227E+02 .484809450E-01-.204693300E-04 .391707780E-08-.279248340E-12    2
-.456695052E+05-.288336460E+02-.321171820E+01 .924083860E-01-.712212230E-04    3
 .295255040E-07-.509148160E-11-.421838470E+05 .417951430E+02                   4
DIPE                    C   6H  14O   1     G    300.00   5000.00 1000.00      1
 .961994133E+01 .527564090E-01-.244349190E-04 .491563770E-08-.360965330E-12    2
-.452985516E+05-.220408754E+02-.207944820E+01 .869029220E-01-.602649600E-04    3
 .209337360E-07-.299614610E-11-.422065600E+05 .378635810E+02                   4
TAME                    C   6H  14O   1     G    300.00   5000.00 1000.00      1
 .102413361E+02 .494717450E-01-.210657300E-04 .406005360E-08-.291140680E-12    2
-.438310029E+05-.257392482E+02-.184725690E+01 .864624650E-01-.624059780E-04    3
 .241227640E-07-.391573010E-11-.407484470E+05 .356637750E+02                   4
C6H5CHO                 C   7H   6O   1     G    300.00   5000.00 1000.00      1
 .151976148E+02 .229544430E-01-.714039470E-05 .736589790E-09 .000000000E+00    2
-.120582935E+05-.546270656E+02-.328352400E+01 .610821620E-01-.279524170E-04    3
 .190203190E-08 .000000000E+00-.599503400E+04 .449259300E+02                   4
C7H8                    C   7H   8          G    300.00   5000.00 1000.00      1
 .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
 .590756417E+03-.294263546E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
 .104046480E-07 .000000000E+00 .469335500E+04 .464073200E+02                   4
C6H5OCH3                C   7H   8O   1     G    300.00   5000.00 1393.00      1
 .203938728E+02 .209088165E-01-.722522263E-05 .112997840E-08-.659097524E-13    2
-.186061425E+05-.862920505E+02-.540888697E+01 .873332441E-01-.739639658E-04    3
 .320208039E-07-.556946955E-11-.102821510E+05 .500696056E+02                   4
CRESOL                  C   7H   8O   1     G    300.00   5000.00 1000.00      1
 .109411883E+02 .359221340E-01-.155859930E-04 .305336930E-08-.221926260E-12    2
-.211837368E+05-.322120090E+02-.410479790E+01 .823735850E-01-.680002460E-04    3
 .287114670E-07-.487123580E-11-.173767210E+05 .440872850E+02                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   5000.00 1000.00      1
 .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
-.176276686E+05-.230348046E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
 .104046480E-07 .000000000E+00-.135250700E+05 .527988700E+02                   4
CH3CH3-C5H6             C   7H  12          G    300.00   5000.00 1000.00      1
 .140192352E+02 .351774100E-01-.121769020E-04 .195853870E-08-.120886390E-12    2
-.562170122E+04-.461295916E+02 .191804150E+01 .620151830E-01-.182958650E-04    3
-.181326460E-07 .113526820E-10-.217165720E+04 .175128710E+02                   4
MCYC6-OQOOH             C   7H  12O   3     G    300.00   5000.00 1380.00      1
 .281047951E+02 .298656134E-01-.103750111E-04 .162883933E-08-.952775107E-13    2
-.587524861E+05-.124642473E+03-.502703972E+01 .104102110E+00-.722526077E-04    3
 .243793077E-07-.320129183E-11-.470307327E+05 .542550536E+02                   4
NC7H14                  C   7H  14          G    300.00   5000.00 1390.00      1
 .206190401E+02 .314852991E-01-.107162057E-04 .165827662E-08-.959911785E-13    2
-.196710875E+05-.822507478E+02-.116533279E+01 .790439806E-01-.496101666E-04    3
 .158569009E-07-.205346433E-11-.117362359E+05 .359871070E+02                   4
MCYC6                   C   7H  14          G    300.00   5000.00 1381.00      1
 .220211359E+02 .332076617E-01-.115857900E-04 .182324838E-08-.106797390E-12    2
-.311719553E+05-.103211614E+03-.890848850E+01 .969226774E-01-.576085500E-04    3
 .148743771E-07-.111357720E-11-.196669630E+05 .657804644E+02                   4
NC7H14O                 C   7H  14O   1     G    300.00   5000.00 1397.00      1
 .231122557E+02 .333659362E-01-.114966228E-04 .179372703E-08-.104427245E-12    2
-.438636425E+05-.993466782E+02-.767475343E+01 .108451023E+00-.827531084E-04    3
 .330380469E-07-.541492429E-11-.334640974E+05 .649157213E+02                   4
NC7H13OOH               C   7H  14O   2     G    300.00   5000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   5000.00 1387.00      1
 .288332529E+02 .320168096E-01-.111508456E-04 .175226159E-08-.102520451E-12    2
-.622309509E+05-.116187714E+03 .152936692E+01 .958173466E-01-.696688520E-04    3
 .269540382E-07-.438728126E-11-.526003608E+05 .306986714E+02                   4
NC7H16                  C   7H  16          G    300.00   5000.00 1000.00      1
 .205103125E+02 .346389640E-01-.107743740E-04 .160399760E-08-.937017530E-13    2
-.326499224E+05-.807081180E+02-.679531340E+00 .810756760E-01-.423279310E-04    3
 .697965770E-08 .837326950E-12-.256907030E+05 .329815600E+02                   4
NC7H15OOH               C   7H  16O   2     G    300.00   5000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
C6H5C2H                 C   8H   6          G    300.00   5000.00 1399.00      1
 .190886756E+02 .170819066E-01-.559393248E-05 .845345947E-09-.482537486E-13    2
 .280711996E+05-.790035627E+02-.377007730E+01 .792380003E-01-.711832819E-04    3
 .324077613E-07-.583009863E-11 .350595597E+05 .405332699E+02                   4
BZFUR                   C   8H   6O   1     G    300.00   5000.00 1000.00      1
 .161267559E+02 .242942790E-01-.882919089E-05 .143722155E-08-.865592465E-13    2
-.574867958E+04-.640564836E+02-.785221476E+00 .396432449E-01 .569751746E-04    3
-.114831806E-06 .519411145E-10 .215748538E+03 .302655928E+02                   4
C6H5C2H3                C   8H   8          G    300.00   5000.00 1000.00      1
 .132118086E+02 .297097690E-01-.100379980E-04 .113030440E-08 .000000000E+00    2
 .112255113E+05-.452965784E+02-.314842000E+01 .733550410E-01-.482478610E-04    3
 .120551240E-07 .000000000E+00 .157685200E+05 .395339300E+02                   4
C6H5C2H5                C   8H  10          G    300.00   5000.00 1000.00      1
 .123967254E+02 .365194120E-01-.128125900E-04 .149467160E-08 .000000000E+00    2
-.304290347E+04-.409211516E+02-.458801200E+01 .813929890E-01-.516055260E-04    3
 .123987680E-07 .000000000E+00 .171000000E+04 .472934500E+02                   4
XYLENE                  C   8H  10          G    300.00   5000.00 1000.00      1
 .104572604E+02 .403200160E-01-.145441770E-04 .173870560E-08 .000000000E+00    2
-.392485555E+04-.316838798E+02-.365621300E+01 .742185790E-01-.400008720E-04    3
 .741031100E-08 .000000000E+00 .307000000E+03 .427477900E+02                   4
UME7                    C   8H  14O   2     G    300.00   5000.00 1386.00      1
 .274195251E+02 .331653074E-01-.112369879E-04 .173174767E-08-.999867016E-13    2
-.597230517E+05-.112624254E+03 .202528941E+01 .898844344E-01-.593620598E-04    3
 .203016355E-07-.286718129E-11-.505953610E+05 .247655861E+02                   4
IC8H16                  C   8H  16          G    300.00   5000.00 1000.00      1
 .159403331E+02 .467083530E-01-.162445520E-04 .262105430E-08-.162114790E-12    2
-.212288474E+05-.575000710E+02-.188446240E+01 .875446570E-01-.337527930E-04    3
-.140196880E-07 .109753600E-10-.160534330E+05 .363096160E+02                   4
IC8H16O                 C   8H  16O   1     G    300.00   5000.00 1400.00      1
 .286870453E+02 .350973257E-01-.120318626E-04 .187165307E-08-.108763411E-12    2
-.489758985E+05-.130519447E+03-.811336944E+01 .120858100E+00-.869108786E-04    3
 .308943900E-07-.431018679E-11-.363657206E+05 .668763983E+02                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   5000.00 1395.00      1
 .329665839E+02 .352889373E-01-.121856584E-04 .190423031E-08-.110989507E-12    2
-.686224367E+05-.138776314E+03 .233137835E+00 .110643301E+00-.779138892E-04    3
 .277663606E-07-.398875833E-11-.571903320E+05 .373387625E+02                   4
IC8H18                  C   8H  18          G    300.00   5000.00 1000.00      1
 .175409498E+02 .499242880E-01-.172020170E-04 .275518900E-08-.169419330E-12    2
-.363533756E+05-.670046390E+02-.203218650E+01 .946845260E-01-.357433050E-04    3
-.165946760E-07 .125346320E-10-.306832730E+05 .359861450E+02                   4
INDENE                  C   9H   8          G    300.00   5000.00 1000.00      1
 .129942100E+02 .345035980E-01-.119473340E-04 .137705200E-08 .000000000E+00    2
 .128398488E+05-.468095535E+02-.565650900E+01 .835992990E-01-.541865810E-04    3
 .131713170E-07 .000000000E+00 .180739000E+05 .501175500E+02                   4
NPBENZ                  C   9H  12          G    300.00   5000.00 1395.00      1
 .234758956E+02 .300348225E-01-.102493106E-04 .158931255E-08-.921475616E-13    2
-.109980792E+05-.102092892E+03-.597461242E+01 .101439137E+00-.768408376E-04    3
 .299742828E-07-.474668103E-11-.108882285E+04 .550543799E+02                   4
TMBENZ                  C   9H  12          G    300.00   5000.00 1383.00      1
 .215885246E+02 .321229102E-01-.110727239E-04 .172825742E-08-.100649304E-12    2
-.136169019E+05-.914142733E+02-.173308850E+01 .786049041E-01-.431048197E-04    3
 .100745302E-07-.585489308E-12-.471446607E+04 .366811038E+02                   4
C7H15COCHO              C   9H  16O   2     G    300.00   5000.00 1387.00      1
 .303225194E+02 .381334789E-01-.128450948E-04 .197085647E-08-.113456990E-12    2
-.668175594E+05-.126355483E+03-.229351926E+00 .108754598E+00-.755330139E-04    3
 .275093508E-07-.415197146E-11-.560981532E+05 .380532571E+02                   4
C10H8                   C  10H   8          G    300.00   5000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
C10H7OH                 C  10H   8O   1     G    300.00   5000.00 1394.00      1
 .262017858E+02 .245473904E-01-.859268465E-05 .135522543E-08-.795056830E-13    2
-.158010339E+05-.119344614E+03-.322687986E+01 .931430619E-01-.687932451E-04    3
 .249753868E-07-.357353464E-11-.568766282E+04 .385570421E+02                   4
C10H10                  C  10H  10          G    300.00   5000.00 2043.00      1
 .196465049E+02 .362867673E-01-.135117921E-04 .222712581E-08-.134868100E-12    2
 .466515480E+04-.883925826E+02-.975555457E+01 .989343734E-01-.593843991E-04    3
 .154882804E-07-.129445409E-11 .148791325E+05 .708155586E+02                   4
TETRALIN                C  10H  12          G    300.00   5000.00 1393.00      1
 .259510150E+02 .311178636E-01-.105072610E-04 .161945272E-08-.935513420E-13    2
-.106963510E+05-.121999608E+03-.103201470E+02 .118533935E+00-.903074920E-04    3
 .343768814E-07-.519161790E-11 .142964373E+04 .715127353E+02                   4
DCYC5                   C  10H  16          G    300.00   5000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
KHDECA                  C  10H  16O   3     G    300.00   5000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
DECALIN                 C  10H  18          G    300.00   5000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
ODECAL                  C  10H  18          G    300.00   5000.00 1383.00      1
 .304308606E+02 .423969327E-01-.145305017E-04 .226051483E-08-.131385276E-12    2
-.274622725E+05-.143201137E+03-.921337866E+01 .127293330E+00-.797537373E-04    3
 .229874961E-07-.227548927E-11-.131010829E+05 .721555536E+02                   4
NC10H20                 C  10H  20          G    300.00   5000.00 1390.00      1
 .306417045E+02 .444757412E-01-.152579717E-04 .237363570E-08-.137907421E-12    2
-.321647483E+05-.129750528E+03-.253770965E+01 .118319727E+00-.776112696E-04    3
 .262647573E-07-.366153318E-11-.202029921E+05 .498650630E+02                   4
NC20MOOH                C  10H  20O   2     G    300.00   5000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   5000.00 1390.00      1
 .373427699E+02 .457774433E-01-.156578702E-04 .243101177E-08-.141046271E-12    2
-.740262240E+05-.156527917E+03 .209018845E+01 .128739739E+00-.918467610E-04    3
 .350282382E-07-.560696315E-11-.617151278E+05 .328016208E+02                   4
NC10H22                 C  10H  22          G    300.00   5000.00 1391.00      1
 .319882239E+02 .477244922E-01-.162276391E-04 .250963259E-08-.145215772E-12    2
-.466392840E+05-.137615344E+03-.208416969E+01 .122535012E+00-.776815739E-04    3
 .249834877E-07-.323548038E-11-.343021863E+05 .471147911E+02                   4
C10H7CHO                C  11H   8O   1     G    300.00   5000.00 1391.00      1
 .276532029E+02 .258287942E-01-.902879433E-05 .142281038E-08-.834251834E-13    2
-.106453206E+05-.124981465E+03-.108527081E+01 .881681978E-01-.575973932E-04    3
 .170999043E-07-.173813923E-11-.356369995E+03 .307785222E+02                   4
C10H7CH3                C  11H  10          G    300.00   5000.00 1394.00      1
 .269623579E+02 .288172394E-01-.100254209E-04 .157466721E-08-.921126923E-13    2
 .586670370E+03-.125206708E+03-.798962224E+01 .117448428E+00-.976360478E-04    3
 .414932114E-07-.710609396E-11 .120022223E+05 .599922187E+02                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   5000.00 1392.00      1
 .281549167E+02 .299236572E-01-.104056239E-04 .163381420E-08-.955470229E-13    2
-.208064399E+05-.126965793E+03-.171335238E+01 .970093442E-01-.665430499E-04    3
 .223717851E-07-.293871610E-11-.102462828E+05 .342637221E+02                   4
UME10                   C  11H  20O   2     G    300.00   5000.00 1384.00      1
 .374112533E+02 .458948435E-01-.156057696E-04 .241315080E-08-.139673864E-12    2
-.736971925E+05-.162545741E+03 .937241013E+00 .126885097E+00-.836053178E-04    3
 .282312118E-07-.390359926E-11-.605539595E+05 .349335674E+02                   4
ETEROMD                 C  11H  20O   3     G    300.00   5000.00 1386.00      1
 .418053606E+02 .443798286E-01-.151698489E-04 .235874245E-08-.137104681E-12    2
-.896960798E+05-.186388223E+03-.869108022E+00 .143689897E+00-.103700029E-03    3
 .384483018E-07-.582555005E-11-.748416098E+05 .429341731E+02                   4
MDKETO                  C  11H  20O   5     G    300.00   5000.00 1391.00      1
 .435827467E+02 .471875465E-01-.155121189E-04 .235632808E-08-.134947249E-12    2
-.114156459E+06-.184940808E+03 .336575533E+01 .147442203E+00-.113482823E-03    3
 .468018272E-07-.796034235E-11-.100759720E+06 .289177372E+02                   4
MD                      C  11H  22O   2     G    300.00   5000.00 1382.00      1
 .393230373E+02 .488368389E-01-.166923510E-04 .259065840E-08-.150309877E-12    2
-.885441006E+05-.173932688E+03 .176901386E+01 .129360919E+00-.808243357E-04    3
 .251676921E-07-.312062272E-11-.747104475E+05 .304352079E+02                   4
C12H8                   C  12H   8          G    300.00   5000.00 1000.00      1
 .213682716E+02 .324830670E-01-.101214580E-04 .104613640E-08 .000000000E+00    2
 .210494631E+05-.924787980E+02-.672892800E+01 .106967800E+00-.747993040E-04    3
 .193364490E-07 .000000000E+00 .288910000E+05 .533672000E+02                   4
DIBZFUR                 C  12H   8O   1     G    300.00   5000.00 1000.00      1
 .238928699E+02 .342239370E-01-.125916314E-04 .206592304E-08-.125089220E-12    2
-.481449779E+04-.107327684E+03-.194754604E+01 .663215475E-01 .555418713E-04    3
-.135401425E-06 .629515620E-10 .401745217E+04 .350605098E+02                   4
BIPHENYL                C  12H  10          G    300.00   5000.00 1000.00      1
 .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
 .115420788E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
 .194042280E-07 .000000000E+00 .198069600E+05 .608493300E+02                   4
DIFENET                 C  12H  10O   1     G    300.00   5000.00 1000.00      1
 .283319364E+02 .317670352E-01-.107447484E-04 .165690065E-08-.957158914E-13    2
-.789446240E+04-.127230446E+03-.865410063E+01 .124988347E+00-.100933530E-03    3
 .413234204E-07-.675938299E-11 .409381103E+04 .686981333E+02                   4
C12H18                  C  12H  18          G    300.00   5000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
C12H22                  C  12H  22          G    300.00   5000.00 1392.00      1
 .362943970E+02 .488870789E-01-.165740715E-04 .255852468E-08-.147868438E-12    2
-.229987583E+05-.159907963E+03-.329755440E+01 .140713318E+00-.978288195E-04    3
 .352594898E-07-.520523450E-11-.920475977E+04 .529246931E+02                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   5000.00 1678.00      1
 .447068212E+02 .522272795E-01-.195350799E-04 .322923457E-08-.195935332E-12    2
-.818914807E+05-.192299360E+03 .877388676E+01 .119113497E+00-.561329021E-04    3
 .677643630E-08 .106366869E-11-.685051188E+05 .572134782E+01                   4
NC12H26                 C  12H  26          G    300.00   5000.00 1391.00      1
 .385099212E+02 .563550048E-01-.191493200E-04 .296024862E-08-.171244150E-12    2
-.548849270E+05-.169785166E+03-.262181594E+01 .147237711E+00-.943970271E-04    3
 .307441268E-07-.403602230E-11-.400654253E+05 .529882396E+02                   4
FLUORENE                C  13H  10          G    300.00   5000.00 1000.00      1
 .231612871E+02 .392128530E-01-.125431510E-04 .133503890E-08 .000000000E+00    2
 .123102892E+05-.103717257E+03-.112092800E+02 .129847800E+00-.907013380E-04    3
 .232288460E-07 .000000000E+00 .219426600E+05 .748524200E+02                   4
C6H5CH2C6H5             C  13H  12          G    300.00   5000.00 1000.00      1
 .185418955E+02 .513343070E-01-.178726910E-04 .207043850E-08 .000000000E+00    2
 .668552054E+04-.690121392E+02-.940899900E+01 .125451300E+00-.822539730E-04    3
 .202856220E-07 .000000000E+00 .144845500E+05 .760677200E+02                   4
ALDINS                  C  13H  20O   1     G    300.00   5000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
U2ME12                  C  13H  22O   2     G    300.00   5000.00 1391.00      1
 .422353117E+02 .524987045E-01-.181261023E-04 .283174793E-08-.165001495E-12    2
-.676968189E+05-.186270028E+03 .679798314E-01 .152530074E+00-.111376081E-03    3
 .435663556E-07-.715842617E-11-.529996239E+05 .399987338E+02                   4
C14H10                  C  14H  10          G    300.00   5000.00 1000.00      1
 .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
 .131224037E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
 .240156710E-07 .000000000E+00 .227649500E+05 .639753600E+02                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   5000.00 1000.00      1
 .183724857E+02 .606470630E-01-.215506390E-04 .254284330E-08 .000000000E+00    2
 .518516081E+04-.659251182E+02-.814781700E+01 .130620600E+00-.819367560E-04    3
 .194757260E-07 .000000000E+00 .126141800E+05 .718458700E+02                   4
C16H10                  C  16H  10          G    300.00   5000.00 1000.00      1
 .290747022E+02 .412337670E-01-.126077060E-04 .127453580E-08 .000000000E+00    2
 .141687238E+05-.136431347E+03-.106811200E+02 .146535400E+00-.103943520E-03    3
 .270645390E-07 .000000000E+00 .252715000E+05 .699617500E+02                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   5000.00 1397.00      1
 .620188250E+02 .682375774E-01-.235322180E-04 .367416933E-08-.214025539E-12    2
-.107194396E+06-.296402060E+03-.700111687E+01 .236135134E+00-.181200158E-03    3
 .715715364E-07-.114883341E-10-.839739066E+05 .717765001E+02                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   5000.00 1854.00      1
 .488264318E+02 .825357366E-01-.292747409E-04 .467245514E-08-.276718037E-12    2
-.942845289E+05-.205583924E+03 .138386904E+01 .198379105E+00-.134722947E-03    3
 .475955890E-07-.691333208E-11-.791319641E+05 .463051187E+02                   4
NC16H34                 C  16H  34          G    300.00   5000.00 1391.00      1
 .515593854E+02 .736064257E-01-.249888737E-04 .386085377E-08-.223263662E-12    2
-.713781425E+05-.234158439E+03-.369111950E+01 .196612966E+00-.127777824E-03    3
 .422323349E-07-.562967041E-11-.515927302E+05 .647080513E+02                   4
IC16H34                 C  16H  34          G    300.00   5000.00 1400.00      1
 .565856523E+02 .692869560E-01-.234931111E-04 .362720220E-08-.209665225E-12    2
-.820366778E+05-.276851694E+03-.107545408E+02 .233995831E+00-.178076331E-03    3
 .696956034E-07-.110282035E-10-.595981394E+05 .818346760E+02                   4
UME16                   C  17H  32O   2     G    300.00   5000.00 1000.00      1
 .333606142E+02 .106719124E+00-.429500189E-04 .790457654E-08-.546125152E-12    2
-.868236054E+05-.126816968E+03 .114310960E+02 .102101194E+00 .102480878E-03    3
-.181385357E-06 .698603588E-10-.778209017E+05 .206428096E+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   5000.00 1000.00      1
 .406345250E+02 .963702350E-01-.332815250E-04 .536978820E-08-.333546480E-12    2
-.105022900E+06-.161181400E+03-.374618910E+01 .216936450E+00-.134184780E-03    3
 .217036750E-07 .800116570E-11-.930412810E+05 .677468110E+02                   4
MPA                     C  17H  34O   2     G    300.00   5000.00 1000.00      1
 .355305296E+02 .109746228E+00-.440981772E-04 .810571172E-08-.559469785E-12    2
-.102923616E+06-.145292419E+03 .117629996E+02 .108027697E+00 .103662595E-03    3
-.187190120E-06 .724616510E-10-.933306777E+05-.643066315E+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   5000.00 1843.00      1
 .597680898E+02 .832144998E-01-.302817533E-04 .491632066E-08-.294624551E-12    2
-.961002787E+05-.258440317E+03-.347354324E+01 .238348931E+00-.171810701E-03    3
 .624560833E-07-.914836595E-11-.760003616E+05 .770024622E+02                   4
MLIN1                   C  19H  32O   2     G    300.00   5000.00 1834.00      1
 .520202170E+02 .871284776E-01-.313984409E-04 .506450961E-08-.302130761E-12    2
-.727531890E+05-.226713941E+03-.298592567E+01 .218746556E+00-.148096154E-03    3
 .511216154E-07-.719451974E-11-.549290521E+05 .662774857E+02                   4
MLINO                   C  19H  34O   2     G    300.00   5000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
MEOLE                   C  19H  36O   2     G    300.00   5000.00 1831.00      1
 .528856562E+02 .948572658E-01-.338668063E-04 .542873444E-08-.322458135E-12    2
-.101075125E+06-.229348639E+03-.267573662E+00 .220639742E+00-.143861659E-03    3
 .481699649E-07-.661786902E-11-.837166223E+05 .542791001E+02                   4
MSTEAKETO               C  19H  36O   5     G    300.00   5000.00 1857.00      1
 .628573476E+02 .927885184E-01-.331648431E-04 .532086973E-08-.316267196E-12    2
-.142644021E+06-.277684268E+03-.711176329E+00 .251338095E+00-.180571731E-03    3
 .664483461E-07-.990089173E-11-.122716422E+06 .585265768E+02                   4
MSTEA                   C  19H  38O   2     G    300.00   5000.00 1000.00      1
 .418174710E+02 .117959830E+00-.465265590E-04 .845319460E-08-.579171090E-12    2
-.110862900E+06-.175601040E+03 .114771030E+02 .131225240E+00 .898738730E-04    3
-.183685190E-06 .722337400E-10-.991500330E+05-.163992920E+01                   4
BIN1B                   C  20H  10          G    300.00   5000.00 1000.00      1
 .228710599E+02 .794839410E-01-.421619700E-04 .106691760E-07-.104891690E-11    2
 .555088663E+05-.100165423E+03-.143921700E+02 .205071170E+00-.201668750E-03    3
 .100637160E-06-.198341200E-10 .644124530E+05 .861129840E+02                   4
BIN1A                   C  20H  16          G    300.00   5000.00 1000.00      1
 .228710599E+02 .794839410E-01-.421619700E-04 .106691760E-07-.104891690E-11    2
 .555088663E+05-.100165423E+03-.143921700E+02 .205071170E+00-.201668750E-03    3
 .100637160E-06-.198341200E-10 .644124530E+05 .861129840E+02                   4
N                       N   1               G    300.00   5000.00 1000.00      1
 .245026778E+01 .106614600E-03-.746533710E-07 .187965200E-10-.102598400E-14    2
 .561160257E+05 .444874779E+01 .250307100E+01-.218001810E-04 .542052910E-07    3
-.564755990E-10 .209990390E-13 .560988900E+05 .416756600E+01                   4
O                       O   1               G    300.00   5000.00 1000.00      1
 .254205876E+01-.275506100E-04-.310280290E-08 .455106700E-11-.436805100E-15    2
 .292307989E+05 .492030884E+01 .294642800E+01-.163816600E-02 .242103100E-05    3
-.160284300E-08 .389069610E-12 .291476400E+05 .296399500E+01                   4
NO3                     O   3N   1          G    300.00   5000.00 1000.00      1
 .712030587E+01 .324622800E-02-.143161340E-05 .279705300E-09-.201300700E-13    2
 .586448126E+04-.121372920E+02 .122107630E+01 .187879700E-01-.134432120E-04    3
 .127460130E-08 .135406010E-11 .747314400E+04 .184020200E+02                   4
H                       H   1               G    300.00   5000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
 .254716200E+05-.460117600E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00 .254716200E+05-.460117600E+00                   4
NH                      H   1N   1          G    300.00   5000.00 1000.00      1
 .276025108E+01 .137534600E-02-.445191400E-06 .769279080E-10-.501759190E-14    2
 .420782748E+05 .585718609E+01 .333975800E+01 .125300900E-02-.349164500E-05    3
 .421881200E-08-.155761800E-11 .418504700E+05 .250718000E+01                   4
NNH                     H   1N   2          G    300.00   5000.00 1000.00      1
 .441534072E+01 .161438800E-02-.163289400E-06-.855984590E-10 .161479110E-13    2
 .278802961E+05 .904297112E+00 .350134400E+01 .205358610E-02 .717040900E-06    3
 .492134780E-09-.967117010E-12 .283334700E+05 .639183800E+01                   4
OH                      H   1O   1          G    300.00   5000.00 1710.00      1
 .285376040E+01 .102994334E-02-.232666477E-06 .193750704E-10-.315759847E-15    2
 .369949720E+04 .578756825E+01 .341896226E+01 .319255801E-03-.308292717E-06    3
 .364407494E-09-.100195479E-12 .345264448E+04 .254433372E+01                   4
HO2                     H   1O   2          G    300.00   5000.00 1000.00      1
 .401721090E+01 .223982013E-02-.633658150E-06 .114246370E-09-.107908535E-13    2
 .111856713E+03 .378510215E+01 .430179801E+01-.474912051E-02 .211582891E-04    3
-.242763894E-07 .929225124E-11 .294808040E+03 .371666245E+01                   4
NH2                     H   2N   1          G    300.00   5000.00 1000.00      1
 .296131091E+01 .293269890E-02-.906360010E-06 .161725700E-09-.120420000E-13    2
 .219197637E+05 .577788090E+01 .343249300E+01 .329953990E-02-.661359990E-05    3
 .859094660E-08-.357204610E-11 .217722700E+05 .309011000E+01                   4
H2NO                    H   2O   1N   1     G    300.00   5000.00 1000.00      1
 .149675000E+01 .889472000E-02-.330837000E-05 .405760000E-09 .000000000E+00    2
 .724825208E+04 .175864616E+02 .267141000E+01 .529823000E-02 .360637000E-06    3
-.841417000E-09 .000000000E+00 .696062900E+04 .116499100E+02                   4
N2H3                    H   3N   2          G    300.00   5000.00 1000.00      1
 .444184100E+01 .721427100E-02-.249568400E-05 .392056500E-09-.229895000E-13    2
 .166422164E+05-.427486304E+00 .317420400E+01 .471590700E-02 .133486700E-04    3
-.191968500E-07 .748756400E-11 .172727000E+05 .755722400E+01                   4
CSOLID                  C   1               G    300.00   5000.00 1000.00      1
 .145569246E+01 .171706380E-02-.697584100E-06 .135283160E-09-.967649050E-14    2
-.695128087E+03-.852568475E+01-.310872070E+00 .440353690E-02 .190394120E-05    3
-.638546970E-08 .298964250E-11-.108650790E+03 .111382950E+01                   4
C                       C   1               G    300.00   5000.00 1000.00      1
 .249266888E+01 .479889284E-04-.724335020E-07 .374291029E-10-.487277893E-14    2
 .854512953E+05 .480150373E+01 .255423955E+01-.321537724E-03 .733792245E-06    3
-.732234889E-09 .266521446E-12 .854438832E+05 .453130848E+01                   4
CN                      C   1N   1          G    300.00   5000.00 1000.00      1
 .372011754E+01 .151835110E-03 .198738110E-06-.379837100E-10 .132823000E-14    2
 .511162563E+05 .288861031E+01 .366320400E+01-.115652890E-02 .216340890E-05    3
 .185420800E-09-.821469520E-12 .512811700E+05 .373901500E+01                   4
NCO                     C   1O   1N   1     G    300.00   5000.00 1000.00      1
 .501204558E+01 .262677300E-02-.110824310E-05 .209385990E-09-.146034700E-13    2
 .173718555E+05-.183007911E+01 .283032000E+01 .887149010E-02-.894563620E-05    3
 .587691810E-08-.190773400E-11 .180054300E+05 .949883200E+01                   4
CH                      C   1H   1          G    300.00   5000.00 1000.00      1
 .219622115E+01 .234038100E-02-.705820130E-06 .900758220E-10-.385504010E-14    2
 .708672121E+05 .917838138E+01 .320020200E+01 .207287490E-02-.513443090E-05    3
 .573388980E-08-.195553300E-11 .704525700E+05 .333158700E+01                   4
HCO                     C   1H   1O   1     G    300.00   5000.00 1000.00      1
 .355727119E+01 .334557190E-02-.133500600E-05 .247057210E-09-.171385000E-13    2
 .391632208E+04 .555229973E+01 .289832900E+01 .619914620E-02-.962308420E-05    3
 .108982500E-07-.457488520E-11 .415992100E+04 .898361500E+01                   4
HCO3                    C   1H   1O   3     G    300.00   5000.00 1368.00      1
 .724073447E+01 .463312951E-02-.163693995E-05 .259706693E-09-.152964699E-13    2
-.187027386E+05-.649534993E+01 .396059309E+01 .106002279E-01-.525713351E-05    3
 .101716726E-08-.287487602E-13-.173599383E+05 .117807483E+02                   4
CH2                     C   1H   2          G    300.00   5000.00 1000.00      1
 .363640757E+01 .193305600E-02-.168701600E-06-.100989900E-09 .180825510E-13    2
 .453413341E+05 .215656196E+01 .376223700E+01 .115981900E-02 .248958490E-06    3
 .880083620E-09-.733243490E-12 .453679000E+05 .171257700E+01                   4
CH2S                    C   1H   2          G    300.00   5000.00 1000.00      1
 .355288641E+01 .206678800E-02-.191411600E-06-.110467300E-09 .202134890E-13    2
 .498497521E+05 .168658499E+01 .397126500E+01-.169908800E-03 .102536900E-05    3
 .249254990E-08-.198126610E-11 .498936700E+05 .575320760E-01                   4
H2CN                    C   1H   2N   1     G    300.00   5000.00 1000.00      1
 .520970151E+01 .296929110E-02-.285558910E-06-.163555000E-09 .304325890E-13    2
 .276771105E+05-.444446452E+01 .285166100E+01 .569523310E-02 .107114000E-05    3
-.162261200E-08-.235110810E-12 .286378200E+05 .899274900E+01                   4
CH3                     C   1H   3          G    300.00   5000.00 1000.00      1
 .284405718E+01 .613797410E-02-.223034500E-05 .378516110E-09-.245215900E-13    2
 .164378004E+05 .545265727E+01 .243044200E+01 .111241000E-01-.168022000E-04    3
 .162182910E-07-.586495220E-11 .164237800E+05 .678979400E+01                   4
CH2OH                   C   1H   3O   1     G    300.00   5000.00 1000.00      1
 .632751914E+01 .360827010E-02-.320154700E-06-.193875000E-09 .350970410E-13    2
-.447450931E+04-.832935988E+01 .286262800E+01 .100152700E-01-.528543520E-06    3
-.513853890E-08 .224604100E-11-.334967800E+04 .103979400E+02                   4
CH3O                    C   1H   3O   1     G    300.00   5000.00 1000.00      1
 .377081447E+01 .787149740E-02-.265638390E-05 .394443090E-09-.211261600E-13    2
 .127818951E+03 .292947482E+01 .210620400E+01 .721659510E-02 .533847200E-05    3
-.737763630E-08 .207561010E-11 .978601200E+03 .131521800E+02                   4
CH3OO                   C   1H   3O   2     G    300.00   5000.00 1385.00      1
 .595784570E+01 .790728626E-02-.268246234E-05 .413891337E-09-.239007330E-13    2
-.378178515E+03-.353671121E+01 .426146906E+01 .100873599E-01-.321506184E-05    3
 .209409267E-09 .418339103E-13 .473129653E+03 .634599067E+01                   4
C2H                     C   2H   1          G    300.00   5000.00 1000.00      1
 .316780603E+01 .475221900E-02-.183787070E-05 .304190250E-09-.177232770E-13    2
 .671210651E+05 .663589763E+01 .288965730E+01 .134099610E-01-.284769500E-04    3
 .294791040E-07-.109331510E-10 .668393930E+05 .622296430E+01                   4
HCCO                    C   2H   1O   1     G    300.00   5000.00 1000.00      1
 .675807437E+01 .200040010E-02-.202760700E-06-.104113200E-09 .196516400E-13    2
 .190151261E+05-.907126528E+01 .504796600E+01 .445347790E-02 .226828210E-06    3
-.148209400E-08 .225074100E-12 .196589100E+05 .481843900E+00                   4
CH2CN                   C   2H   2N   1     G    300.00   5000.00 1000.00      1
 .460581482E+01 .944851600E-02-.471163290E-05 .113899570E-08-.108289420E-12    2
 .291714861E+05 .100843943E+01 .252967240E+01 .181141380E-01-.189605750E-04    3
 .119445830E-07-.325441420E-11 .295922930E+05 .109934410E+02                   4
C2H3                    C   2H   3          G    300.00   5000.00 1000.00      1
 .593346697E+01 .401774510E-02-.396673900E-06-.144126700E-09 .237864300E-13    2
 .318543468E+05-.853030497E+01 .245927600E+01 .737147590E-02 .210987200E-05    3
-.132164200E-08-.118478400E-11 .333522500E+05 .115562000E+02                   4
CH3CO                   C   2H   3O   1     G    300.00   5000.00 1000.00      1
 .561230883E+01 .844988600E-02-.285414690E-05 .423837600E-09-.226840300E-13    2
-.518788372E+04-.327515155E+01 .312527800E+01 .977822020E-02 .452144790E-05    3
-.900946160E-08 .319371700E-11-.410850700E+04 .112288500E+02                   4
CH2CHO                  C   2H   3O   1     G    300.00   5000.00 1500.00      1
 .971005743E+01 .385496600E-02-.467782500E-06-.150517900E-09 .294142800E-13    2
-.269248263E+04-.281056408E+02 .280220500E+00 .274031100E-01-.255468300E-04    3
 .130667900E-07-.275042500E-11 .668264800E+03 .223973100E+02                   4
CH3OCO                  C   2H   3O   2     G    300.00   5000.00 1601.00      1
 .973659803E+01 .742432713E-02-.265641779E-05 .425031143E-09-.251824924E-13    2
-.235512450E+05-.237360013E+02 .416215406E+01 .138037511E-01-.308486109E-06    3
-.456430814E-08 .146909632E-11-.209627030E+05 .854235619E+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   5000.00 1000.00      1
 .102188027E+02 .888408630E-02-.222887620E-05 .166265570E-09 .000000000E+00    2
-.256023886E+05-.219354293E+02 .384065500E+01 .218595100E-01-.904528040E-05    3
 .385393800E-09 .000000000E+00-.234946000E+05 .124829900E+02                   4
C2H5                    C   2H   5          G    300.00   5000.00 1000.00      1
 .719047846E+01 .648407680E-02-.642806410E-06-.234787910E-09 .388087690E-13    2
 .106745471E+05-.147808755E+02 .269070100E+01 .871913320E-02 .441983820E-05    3
 .933870310E-09-.392777300E-11 .128704000E+05 .121382000E+02                   4
CH3CHOH                 C   2H   5O   1     G    300.00   5000.00 1553.00      1
 .726570301E+01 .109588926E-01-.363662803E-05 .553659830E-09-.317012322E-13    2
-.864371441E+04-.106822851E+02 .183974631E+01 .187789371E-01-.460544253E-05    3
-.213116990E-08 .943772653E-12-.629595195E+04 .201446141E+02                   4
C2H4OH                  C   2H   5O   1     G    300.00   5000.00 1391.00      1
 .752244726E+01 .110492715E-01-.372576465E-05 .572827397E-09-.330061759E-13    2
-.729337464E+04-.124960750E+02 .117714711E+01 .248115685E-01-.150299503E-04    3
 .479006785E-08-.640994211E-12-.495369043E+04 .220081586E+02                   4
CH3OCH2                 C   2H   5O   1     G    300.00   5000.00 1376.00      1
 .817131769E+01 .110086181E-01-.382352277E-05 .599637202E-09-.350317513E-13    2
-.291606126E+04-.178646468E+02 .291327415E+01 .203364659E-01-.959712342E-05    3
 .207478525E-08-.171343362E-12-.685171134E+03 .116066817E+02                   4
C2H5OO                  C   2H   5O   2     G    300.00   5000.00 1388.00      1
 .951115499E+01 .122676900E-01-.422364452E-05 .658474989E-09-.383095208E-13    2
-.676067578E+04-.223427083E+02 .177950508E+01 .304938087E-01-.216376209E-04    3
 .868906296E-08-.151788464E-11-.399101974E+04 .192919501E+02                   4
C2-QOOH                 C   2H   5O   2     G    300.00   5000.00 1396.00      1
 .116258666E+02 .100826346E-01-.347934362E-05 .543394220E-09-.316569294E-13    2
-.910568267E+03-.318522902E+02 .813237801E+00 .390063400E-01-.340643855E-04    3
 .155066226E-07-.284069840E-11 .250785787E+04 .249684459E+02                   4
DME-QOOH                C   2H   5O   3     G    300.00   5000.00 1367.00      1
 .140894827E+02 .105710448E-01-.375281006E-05 .597314407E-09-.352604582E-13    2
-.191406716E+05-.429268872E+02 .543520255E+01 .272005914E-01-.150210893E-04    3
 .370396290E-08-.309396378E-12-.157034464E+05 .495012674E+01                   4
DME-OO                  C   2H   5O   3     G    300.00   5000.00 1359.00      1
 .120501213E+02 .123072703E-01-.435221905E-05 .690896352E-09-.407091104E-13    2
-.227977573E+05-.323415629E+02 .515628105E+01 .216783339E-01-.561847228E-05    3
-.192807296E-08 .859447044E-12-.196244836E+05 .725163812E+01                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   5000.00 1387.00      1
 .145471032E+02 .123393823E-01-.427259469E-05 .668763337E-09-.390196721E-13    2
-.196338761E+05-.408784236E+02 .590031872E+01 .305658528E-01-.185905950E-04    3
 .567871605E-08-.702799577E-12-.163916571E+05 .633051038E+01                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   5000.00 1382.00      1
 .146274659E+02 .163794767E-01-.563311171E-05 .877481381E-09-.510186598E-13    2
-.370029335E+05-.399555488E+02 .771229157E+01 .301140957E-01-.165996092E-04    3
 .533577253E-08-.842885930E-12-.341808026E+05-.165902348E+01                   4
C3H3                    C   3H   3          G    300.00   5000.00 1000.00      1
 .883104772E+01 .435719410E-02-.410906610E-06-.236872300E-09 .437652000E-13    2
 .384741917E+05-.217791939E+02 .475419900E+01 .110802800E-01 .279332310E-06    3
-.547921220E-08 .194962900E-11 .398888300E+05 .585454700E+00                   4
CH2CHCH2                C   3H   5          G    300.00   5000.00 1000.00      1
 .846871473E+01 .110576240E-01-.329817360E-05 .323385870E-09 .000000000E+00    2
 .160467269E+05-.206696057E+02 .227648600E+01 .198556410E-01 .112384200E-05    3
-.101457600E-07 .344134200E-11 .182949600E+05 .137251500E+02                   4
CH2CCH3                 C   3H   5          G    300.00   5000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
CHCHCH3                 C   3H   5          G    300.00   5000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
C2H4CHO                 C   3H   5O   1     G    300.00   5000.00 1683.00      1
 .813285396E+01 .137651720E-01-.486366739E-05 .775334875E-09-.459117207E-13    2
-.292071282E+04-.132464943E+02 .324839539E+01 .209600531E-01-.607665825E-05    3
-.115341896E-08 .627874009E-12-.913395491E+03 .143591941E+02                   4
CH3COCH2                C   3H   5O   1     G    300.00   5000.00 1391.00      1
 .102303674E+02 .116494161E-01-.401005537E-05 .625205246E-09-.363784362E-13    2
-.844376284E+04-.279195044E+02 .180339187E+01 .301407085E-01-.193505552E-04    3
 .638199034E-08-.866103180E-12-.537233261E+04 .178046408E+02                   4
C3H5OO                  C   3H   5O   2     G    300.00   5000.00 1375.00      1
 .120289627E+02 .126220050E-01-.443107280E-05 .699998849E-09-.411059161E-13    2
 .440592543E+04-.346276747E+02 .316765415E+01 .300862111E-01-.169786280E-04    3
 .462955698E-08-.501220245E-12 .789477349E+04 .142601307E+02                   4
IC3H7                   C   3H   7          G    300.00   5000.00 1000.00      1
 .736341098E+01 .171331520E-01-.582028000E-05 .658834320E-09 .000000000E+00    2
 .604684608E+04-.148406654E+02 .171329900E+01 .254261610E-01 .158080800E-05    3
-.182128610E-07 .882771030E-11 .803580600E+04 .162790100E+02                   4
NC3H7                   C   3H   7          G    300.00   5000.00 1000.00      1
 .722715260E+01 .172648710E-01-.588880490E-05 .669183600E-09 .000000000E+00    2
 .782835831E+04-.127978858E+02 .192253600E+01 .247892700E-01 .181024900E-05    3
-.178326490E-07 .858299630E-11 .971328300E+04 .164927100E+02                   4
NC3H7O                  C   3H   7O   1     G    300.00   5000.00 1390.00      1
 .107032043E+02 .160908541E-01-.548805425E-05 .850429828E-09-.492755368E-13    2
-.101405419E+05-.313058764E+02-.595838475E+00 .410450833E-01-.263340323E-04    3
 .872638287E-08-.119115039E-11-.604569631E+04 .299328965E+02                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   5000.00 1392.00      1
 .106573810E+02 .155684549E-01-.527663821E-05 .814099260E-09-.470228616E-13    2
-.112728087E+05-.272448749E+02 .975268381E+00 .369225253E-01-.232066980E-04    3
 .768472523E-08-.106762046E-11-.774554528E+04 .252661698E+02                   4
C3H6OH                  C   3H   7O   1     G    300.00   5000.00 1674.00      1
 .931264447E+01 .167567524E-01-.575483066E-05 .900436230E-09-.526465859E-13    2
-.119156359E+05-.195563575E+02 .120238342E+01 .330977268E-01-.164088500E-04    3
 .319283457E-08-.708290455E-13-.902825324E+04 .246699783E+02                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   5000.00 1388.00      1
 .110944203E+02 .153549108E-01-.523574640E-05 .810964124E-09-.469665855E-13    2
-.134769536E+05-.307070215E+02 .584672920E+00 .407370189E-01-.294865043E-04    3
 .116950656E-07-.196228356E-11-.984929391E+04 .255429190E+02                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   5000.00 1674.00      1
 .931287816E+01 .167579212E-01-.575555480E-05 .900584362E-09-.526566836E-13    2
-.119163093E+05-.195564662E+02 .120494302E+01 .330857885E-01-.163893637E-04    3
 .318103918E-08-.684229288E-13-.902896295E+04 .246601603E+02                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   5000.00 1386.00      1
 .110500439E+02 .152562747E-01-.517257413E-05 .798146428E-09-.461030406E-13    2
-.142779432E+05-.312276095E+02 .149130595E+01 .376502110E-01-.258507542E-04    3
 .978662277E-08-.158835656E-11-.109017244E+05 .201908977E+02                   4
CH3COHCH3               C   3H   7O   1     G    300.00   5000.00 1388.00      1
 .115026438E+02 .149881248E-01-.510421075E-05 .789864272E-09-.457135659E-13    2
-.164821894E+05-.347655748E+02 .118802517E+01 .410410262E-01-.314650841E-04    3
 .133514692E-07-.237788249E-11-.130177234E+05 .200655998E+02                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   5000.00 1386.00      1
 .114171877E+02 .153513978E-01-.529698955E-05 .827233821E-09-.481919070E-13    2
-.102618580E+05-.351878119E+02 .408331131E+00 .386748099E-01-.236531335E-04    3
 .722163698E-08-.882900722E-12-.615994143E+04 .248520294E+02                   4
NC3H7OO                 C   3H   7O   2     G    300.00   5000.00 1388.00      1
 .127230991E+02 .167336808E-01-.575943184E-05 .897769493E-09-.522275065E-13    2
-.108816595E+05-.381965321E+02 .156301709E+01 .426192697E-01-.296615075E-04    3
 .114187326E-07-.189894471E-11-.688086375E+04 .219842933E+02                   4
NC3-QOOH                C   3H   7O   2     G    300.00   5000.00 1374.00      1
 .146139980E+02 .143723015E-01-.488635144E-05 .756519620E-09-.438364992E-13    2
-.646101457E+04-.457478245E+02 .191005011E+01 .411666833E-01-.251630217E-04    3
 .711856873E-08-.698838732E-12-.179305093E+04 .234514457E+02                   4
IC3H7OO                 C   3H   7O   2     G    300.00   5000.00 1392.00      1
 .132610651E+02 .162501084E-01-.558631798E-05 .870057473E-09-.505849469E-13    2
-.131937089E+05-.421023499E+02 .103495454E+01 .469942369E-01-.366525520E-04    3
 .157084173E-07-.281956117E-11-.906344820E+04 .229566921E+02                   4
IC3-QOOH                C   3H   7O   2     G    300.00   5000.00 1399.00      1
 .155030898E+02 .139802008E-01-.481811216E-05 .751835399E-09-.437743118E-13    2
-.741643030E+04-.523911482E+02-.184042862E+00 .564670638E-01-.501611253E-04    3
 .230526863E-07-.423866481E-11-.252333896E+04 .298354826E+02                   4
C3H6OHOO                C   3H   7O   3     G    300.00   5000.00 1394.00      1
 .144153388E+02 .176838629E-01-.605016347E-05 .939176426E-09-.544740069E-13    2
-.311104412E+05-.431485877E+02 .184066306E+01 .504311170E-01-.405822327E-04    3
 .181227136E-07-.336967699E-11-.269499345E+05 .234072195E+02                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   5000.00 1391.00      1
 .191234208E+02 .158457151E-01-.552231946E-05 .868162288E-09-.508094203E-13    2
-.255253957E+05-.661419362E+02 .175906535E+01 .624712381E-01-.554930416E-04    3
 .257973727E-07-.483190839E-11-.200009572E+05 .251348546E+02                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   5000.00 1388.00      1
 .185146106E+02 .164157074E-01-.573085844E-05 .901975314E-09-.528299084E-13    2
-.231819444E+05-.618247164E+02 .254387733E+01 .570847379E-01-.472164204E-04    3
 .208289492E-07-.378162942E-11-.178600410E+05 .229447574E+02                   4
C4H3                    C   4H   3          G    300.00   5000.00 1000.00      1
 .107527376E+02 .538115300E-02-.554963720E-06-.305226590E-09 .576173970E-13    2
 .612141980E+05-.297302533E+02 .415388100E+01 .172628700E-01-.238937390E-06    3
-.101870000E-07 .434050410E-11 .633807200E+05 .603650600E+01                   4
C4H5                    C   4H   5          G    300.00   5000.00 1000.00      1
 .128659744E+02 .794336940E-02-.862646570E-06-.465563500E-09 .895113110E-13    2
 .378355213E+05-.418250446E+02 .299524000E+01 .228845610E-01 .197547090E-05    3
-.114824500E-07 .319782310E-11 .414221800E+05 .128945400E+02                   4
IC4H7                   C   4H   7          G    300.00   5000.00 1000.00      1
 .616543300E+01 .257842760E-01-.936521250E-05 .112618500E-08 .000000000E+00    2
 .114713700E+05-.676561500E+01 .476952000E+01 .167724920E-01 .213011010E-04    3
-.275874430E-07 .845501100E-11 .126384700E+05 .401309300E+01                   4
SC4H7                   C   4H   7          G    300.00   5000.00 1000.00      1
 .714879043E+01 .219663880E-01-.774471300E-05 .907477370E-09 .000000000E+00    2
 .124589843E+05-.117547735E+02-.442598200E+00 .422160100E-01-.254697900E-04    3
 .597432100E-08 .000000000E+00 .145672100E+05 .276086500E+02                   4
CH2C3H5                 C   4H   7          G    300.00   5000.00 1000.00      1
 .664945270E+01 .226232110E-01-.806420670E-05 .954149200E-09 .000000000E+00    2
 .206794519E+05-.786429084E+01 .283048200E+00 .386777000E-01-.210739710E-04    3
 .427582900E-08 .000000000E+00 .225247800E+05 .254564400E+02                   4
RMP3                    C   4H   7O   2     G    300.00   5000.00 1376.00      1
 .154260382E+02 .169789201E-01-.593961909E-05 .936106835E-09-.548809672E-13    2
-.343012110E+05-.525677530E+02 .406577480E+01 .388324925E-01-.208048750E-04    3
 .506251249E-08-.421741752E-12-.297848227E+05 .102796868E+02                   4
NC4H9S                  C   4H   9          G    300.00   5000.00 1000.00      1
 .182440000E+01 .354350280E-01-.136901980E-04 .172985780E-08 .000000000E+00    2
 .521137543E+04 .190721830E+02 .882678800E+00 .419813690E-01-.239577090E-04    3
 .639274900E-08 .000000000E+00 .513670700E+04 .226104800E+02                   4
NC4H9P                  C   4H   9          G    300.00   5000.00 1000.00      1
 .285927140E+01 .339093470E-01-.129634890E-04 .162487360E-08 .000000000E+00    2
 .644131902E+04 .136765387E+02 .361027200E+00 .446560900E-01-.269622400E-04    3
 .737512580E-08 .000000000E+00 .679487900E+04 .252696800E+02                   4
IC4H9T                  C   4H   9          G    300.00   5000.00 1000.00      1
 .678309830E+01 .275756420E-01-.999251920E-05 .119923980E-08 .000000000E+00    2
 .130943964E+04-.110379681E+02-.668177200E+00 .478197410E-01-.281268890E-04    3
 .654078610E-08 .000000000E+00 .334806900E+04 .274761900E+02                   4
IC4H9P                  C   4H   9          G    300.00   5000.00 1000.00      1
 .672898190E+01 .277240280E-01-.100574610E-04 .120817530E-08 .000000000E+00    2
 .390175463E+04-.921990655E+01-.514098700E+00 .469939600E-01-.268680800E-04    3
 .599194290E-08 .000000000E+00 .591746700E+04 .283543100E+02                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   5000.00 1389.00      1
 .146211284E+02 .192812832E-01-.662005863E-05 .103030580E-08-.598746774E-13    2
-.185860609E+05-.491894138E+02 .151231967E+01 .485940354E-01-.319829373E-04    3
 .112440534E-07-.168373464E-11-.138241933E+05 .218089522E+02                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   5000.00 1390.00      1
 .151619233E+02 .189741815E-01-.654734215E-05 .102237774E-08-.595503510E-13    2
-.208549516E+05-.532957109E+02 .108860217E+01 .524153990E-01-.380997951E-04    3
 .151074363E-07-.254404184E-11-.159195374E+05 .222613243E+02                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   5000.00 1422.00      1
 .140854789E+02 .197806925E-01-.671026390E-05 .103599950E-08-.598718336E-13    2
-.165129917E+05-.457671006E+02-.566170728E-01 .523981203E-01-.356379876E-04    3
 .128198684E-07-.192264202E-11-.115334457E+05 .303769293E+02                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   5000.00 1673.00      1
 .145354872E+02 .193544788E-01-.655352544E-05 .101052180E-08-.583473661E-13    2
-.195307842E+05-.500528678E+02 .524328525E+00 .528985884E-01-.379651080E-04    3
 .147054933E-07-.239054621E-11-.147012758E+05 .249822692E+02                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   5000.00 1388.00      1
 .142154423E+02 .196229836E-01-.673796562E-05 .104876785E-08-.609536943E-13    2
-.155756339E+05-.451352578E+02 .916505889E+00 .482692226E-01-.299841815E-04    3
 .956515610E-08-.126002465E-11-.106572242E+05 .272437766E+02                   4
CH3CHCH2OCH3            C   4H   9O   1     G    300.00   5000.00 1422.00      1
 .148239632E+02 .195938055E-01-.674334212E-05 .105133556E-08-.611769464E-13    2
-.154937986E+05-.535942326E+02-.581327100E+00 .539666459E-01-.358338761E-04    3
 .122179671E-07-.171024843E-11-.995421675E+04 .297619860E+02                   4
RTC4H8OH                C   4H   9O   1     G    300.00   5000.00 1395.00      1
 .146782533E+02 .193935063E-01-.660052048E-05 .102120044E-08-.590998119E-13    2
-.199408575E+05-.505292168E+02-.836665970E-01 .558040633E-01-.420184309E-04    3
 .171111519E-07-.290735214E-11-.149499995E+05 .281627857E+02                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   5000.00 2017.00      1
 .125195208E+02 .211308942E-01-.735078190E-05 .116027279E-08-.682567448E-13    2
-.159698333E+05-.352643597E+02 .927266773E+00 .453885784E-01-.244944451E-04    3
 .574420616E-08-.382704524E-12-.119074306E+05 .276532069E+02                   4
CH3CH2CHOCH3            C   4H   9O   1     G    300.00   5000.00 1382.00      1
 .157118766E+02 .189436692E-01-.663728010E-05 .104718616E-08-.614402720E-13    2
-.169625442E+05-.584079611E+02-.123566480E+00 .537328693E-01-.359804830E-04    3
 .125064763E-07-.182873667E-11-.111514942E+05 .275750096E+02                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   5000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   5000.00 1387.00      1
 .142049192E+02 .195897318E-01-.671801693E-05 .104483881E-08-.606940644E-13    2
-.190416934E+05-.463876157E+02 .933300006E+00 .472805232E-01-.278316313E-04    3
 .797039080E-08-.870532264E-12-.140666468E+05 .261224696E+02                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   5000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   5000.00 1682.00      1
 .125605997E+02 .210637488E-01-.715019648E-05 .110439262E-08-.638428695E-13    2
-.183183621E+05-.368996627E+02 .329612707E+01 .347649647E-01-.102505618E-04    3
-.204641931E-08 .118879408E-11-.142607619E+05 .157499123E+02                   4
RTC4H9O                 C   4H   9O   1     G    300.00   5000.00 1391.00      1
 .154820006E+02 .191120896E-01-.659337031E-05 .102954283E-08-.599712426E-13    2
-.189474281E+05-.587209701E+02-.652960434E+00 .575360662E-01-.423660204E-04    3
 .165461682E-07-.269335532E-11-.133634774E+05 .277645681E+02                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   5000.00 2017.00      1
 .125195208E+02 .211308942E-01-.735078190E-05 .116027279E-08-.682567448E-13    2
-.159698333E+05-.352643597E+02 .927266773E+00 .453885784E-01-.244944451E-04    3
 .574420616E-08-.382704524E-12-.119074306E+05 .276532069E+02                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   5000.00 1383.00      1
 .150639724E+02 .192754979E-01-.670246160E-05 .105215438E-08-.615166356E-13    2
-.145981078E+05-.535775104E+02 .266423313E+00 .503656318E-01-.308368147E-04    3
 .928122753E-08-.110203449E-11-.905887861E+04 .272172881E+02                   4
NC4-QOOH                C   4H   9O   2     G    300.00   5000.00 1391.00      1
 .182943014E+02 .184250091E-01-.627217889E-05 .971379578E-09-.562825607E-13    2
-.128564704E+05-.650917535E+02 .986162058E+00 .585630676E-01-.416710545E-04    3
 .151223447E-07-.222454695E-11-.684048054E+04 .279289603E+02                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   5000.00 1397.00      1
 .188631296E+02 .183239932E-01-.631233086E-05 .984688082E-09-.573186521E-13    2
-.138981290E+05-.708829284E+02-.425033602E+00 .698121411E-01-.606175877E-04    3
 .274812344E-07-.501908797E-11-.779203954E+04 .305104370E+02                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   5000.00 1396.00      1
 .181457399E+02 .188972595E-01-.650258715E-05 .101363925E-08-.589752496E-13    2
-.103249571E+05-.654833345E+02-.253900783E+00 .658110437E-01-.535280232E-04    3
 .228723790E-07-.398637599E-11-.429699727E+04 .319918975E+02                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   5000.00 1391.00      1
 .160321835E+02 .211162441E-01-.726598082E-05 .113244436E-08-.658740064E-13    2
-.161760498E+05-.559920048E+02 .591660961E+00 .579744782E-01-.422019324E-04    3
 .167841571E-07-.283252682E-11-.107815683E+05 .268393730E+02                   4
NC4H9-OO                C   4H   9O   2     G    300.00   5000.00 1392.00      1
 .164199470E+02 .207668293E-01-.714061871E-05 .111233445E-08-.646799300E-13    2
-.172909027E+05-.576444825E+02 .859225542E+00 .589774363E-01-.445935184E-04    3
 .184502497E-07-.321329944E-11-.119598721E+05 .254554544E+02                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   5000.00 1392.00      1
 .167547908E+02 .205266172E-01-.706765238E-05 .110199004E-08-.641203511E-13    2
-.197490954E+05-.625129056E+02 .429458545E+00 .619305024E-01-.492178248E-04    3
 .213391061E-07-.385156685E-11-.142778206E+05 .242205126E+02                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   5000.00 1393.00      1
 .231119306E+02 .196469811E-01-.682730172E-05 .107124796E-08-.626109519E-13    2
-.320261199E+05-.872192509E+02 .109604492E+01 .794472856E-01-.714221316E-04    3
 .334124791E-07-.626730135E-11-.251118713E+05 .282288973E+02                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   5000.00 1391.00      1
 .225796674E+02 .201772761E-01-.702773819E-05 .110438266E-08-.646157968E-13    2
-.320684788E+05-.852469773E+02 .152317721E+01 .757827720E-01-.656981278E-04    3
 .300159936E-07-.556277284E-11-.252715176E+05 .257762885E+02                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   5000.00 1390.00      1
 .218612263E+02 .207812365E-01-.723484570E-05 .113659545E-08-.664871920E-13    2
-.284979533E+05-.798472350E+02 .156900216E+01 .724191880E-01-.596183448E-04    3
 .260680737E-07-.468228506E-11-.217597632E+05 .278260039E+02                   4
CYC5H5                  C   5H   5          G    300.00   5000.00 1000.00      1
 .421464919E+01 .271834728E-01-.133173209E-04 .308980119E-08-.277879873E-12    2
 .288952416E+05-.305999781E-01-.737844042E+01 .972391818E-01-.169579138E-03    3
 .151818667E-06-.512075479E-10 .305514662E+05 .512829539E+02                   4
C5H5O                   C   5H   5O   1     G    300.00   5000.00 1395.00      1
 .149072105E+02 .136369619E-01-.470762207E-05 .736028654E-09-.429314124E-13    2
 .143724130E+05-.569296345E+02-.414628450E+01 .623584874E-01-.528374678E-04    3
 .224628793E-07-.380136191E-11 .204992627E+05 .437921058E+02                   4
C5H7                    C   5H   7          G    300.00   5000.00 1000.00      1
 .671323690E+01 .274278890E-01-.994311090E-05 .119373240E-08 .000000000E+00    2
 .235116384E+05-.112735252E+02 .759315300E+00 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .251686000E+05 .196131100E+02                   4
CYC5H7                  C   5H   7          G    300.00   5000.00 1416.00      1
 .136844595E+02 .164476117E-01-.550085934E-05 .841117914E-09-.482809780E-13    2
 .196899733E+05-.611528610E+02-.236726157E+01 .584423190E-01-.478622325E-04    3
 .202710415E-07-.344123135E-11 .247432754E+05 .233377340E+02                   4
RMCROTA                 C   5H   7O   2     G    300.00   5000.00 1000.00      1
 .151681730E+02 .178142000E-01-.496258460E-05 .688767770E-09-.386765100E-13    2
-.320532540E+05-.462913590E+02-.242828070E+00 .630479530E-01-.556979940E-04    3
 .265678430E-07-.501508770E-11-.278218120E+05 .329157640E+02                   4
NC5H9                   C   5H   9          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-4                 C   5H   9          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-3                 C   5H   9          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-5                 C   5H   9          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
C5EN-QOOH-54            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO-5               C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C5EN-QOOH-35            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-QOOH-45            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO-3               C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C5EN-QOOH-53            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO-4               C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C5EN-QOOH-43            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
RMBX                    C   5H   9O   2     G    300.00   5000.00 1382.00      1
 .193382201E+02 .209401493E-01-.732209753E-05 .115371679E-08-.676297088E-13    2
-.412852468E+05-.755834444E+02 .231680806E+01 .569247905E-01-.356059275E-04    3
 .110212330E-07-.136558032E-11-.349304634E+05 .172843303E+02                   4
C5EN-QOOH-34            C   5H   9O   2     G    300.00   5000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OOQOOH-43          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-45          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-53          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-54          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
RMBOOX                  C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-34          C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
QMBOOX                  C   5H   9O   4     G    300.00   5000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
ZMBOOX                  C   5H   9O   6     G    300.00   5000.00 1000.00      1
 .261471200E+02 .215283560E-01-.581135510E-05 .785452200E-09-.431572980E-13    2
-.689643590E+05-.913329620E+02 .443715430E+01 .699071290E-01-.165602940E-04    3
-.356586160E-07 .205531550E-10-.628690510E+05 .226288070E+02                   4
NC5H11                  C   5H  11          G    300.00   5000.00 1384.00      1
 .131340658E+02 .260923466E-01-.897731137E-05 .139920325E-08-.813970860E-13    2
-.427735231E+04-.434455998E+02-.304386354E+01 .581995422E-01-.316090839E-04    3
 .790004927E-08-.665198232E-12 .199185425E+04 .455946950E+02                   4
NEOC5H11                C   5H  11          G    300.00   5000.00 1396.00      1
 .166235914E+02 .227037884E-01-.771624835E-05 .119289853E-08-.690060600E-13    2
-.396429146E+04-.644693953E+02-.158140132E+01 .657175067E-01-.468120314E-04    3
 .174732793E-07-.268709925E-11 .230933742E+04 .331296742E+02                   4
RMTBE                   C   5H  11O   1     G    300.00   5000.00 1386.00      1
 .191923401E+02 .226496418E-01-.770522799E-05 .119249279E-08-.690514122E-13    2
-.223486482E+05-.717004889E+02-.284403552E+00 .706092470E-01-.543641242E-04    3
 .224557925E-07-.385680161E-11-.157511970E+05 .321647207E+02                   4
C5H10-OH                C   5H  11O   1     G    300.00   5000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
NC5H12OO                C   5H  11O   2     G    300.00   5000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   5000.00 1396.00      1
 .202154849E+02 .245786365E-01-.841704919E-05 .130775217E-08-.759095109E-13    2
-.224777899E+05-.796085899E+02 .730403748E+00 .705036948E-01-.502866599E-04    3
 .189083885E-07-.294948183E-11-.157211898E+05 .249439750E+02                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   5000.00 1396.00      1
 .218550366E+02 .228989820E-01-.786956915E-05 .122572909E-08-.712760383E-13    2
-.164801773E+05-.857429310E+02 .115441893E+01 .724266160E-01-.535668095E-04    3
 .205704339E-07-.323425526E-11-.941504872E+04 .250054329E+02                   4
NC5-QOOH                C   5H  11O   2     G    300.00   5000.00 1396.00      1
 .220245928E+02 .228314385E-01-.786198359E-05 .122609365E-08-.713571493E-13    2
-.179960313E+05-.864387261E+02-.607426660E+00 .818016374E-01-.685494236E-04    3
 .302071532E-07-.540750321E-11-.106868081E+05 .330450153E+02                   4
C5H10-OHOO              C   5H  11O   3     G    300.00   5000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   5000.00 1401.00      1
 .214971173E+02 .259064341E-01-.848605930E-05 .127921441E-08-.726936886E-13    2
-.312441531E+05-.765479844E+02 .134883146E+01 .795292274E-01-.643595941E-04    3
 .280404405E-07-.497823206E-11-.249060790E+05 .293286141E+02                   4
MTBE-OO                 C   5H  11O   3     G    300.00   5000.00 1386.00      1
 .219476262E+02 .253064866E-01-.877948807E-05 .137597948E-08-.803553517E-13    2
-.383949561E+05-.811182382E+02 .226233362E+01 .712292692E-01-.511734982E-04    3
 .199100134E-07-.329751069E-11-.314029562E+05 .248780910E+02                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   5000.00 1392.00      1
 .248490803E+02 .252599638E-01-.873651764E-05 .136662251E-08-.797082603E-13    2
-.350133010E+05-.961825156E+02 .265748524E+01 .758789336E-01-.526594216E-04    3
 .186692316E-07-.269820831E-11-.271776626E+05 .234450387E+02                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   5000.00 1391.00      1
 .257270270E+02 .247172056E-01-.859292907E-05 .134865114E-08-.788382618E-13    2
-.361631686E+05-.100728579E+03 .135798731E+01 .877212925E-01-.735867140E-04    3
 .327395450E-07-.595540146E-11-.281695250E+05 .282261555E+02                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   5000.00 1391.00      1
 .264681284E+02 .261757287E-01-.899393547E-05 .140058534E-08-.814301239E-13    2
-.504985383E+05-.992053288E+02 .454595241E+01 .801871705E-01-.616423289E-04    3
 .254521416E-07-.437448229E-11-.430642384E+05 .177072264E+02                   4
C6H3                    C   6H   3          G    300.00   5000.00 1000.00      1
 .127611810E+02 .103855730E-01-.347919200E-05 .510973300E-09-.269096500E-13    2
 .747770600E+05-.389174500E+02 .500708900E+01 .269285100E-01-.591986500E-05    3
-.152723350E-07 .940831000E-11 .771320000E+05 .222562100E+01                   4
LC6H5                   C   6H   5          G    300.00   5000.00 1000.00      1
 .134117680E+02 .147202210E-01-.508177050E-05 .798863540E-09-.469508440E-13    2
 .585037160E+05-.416520320E+02 .779297070E+00 .543721260E-01-.478738140E-04    3
 .161871640E-07 .337357440E-12 .616503120E+05 .221285920E+02                   4
C6H5                    C   6H   5          G    300.00   5000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
C6H5O                   C   6H   5O   1     G    300.00   5000.00 1000.00      1
 .137221720E+02 .174688771E-01-.635504520E-05 .103492308E-08-.623410504E-13    2
 .287274751E+03-.488181680E+02-.466204455E+00 .413443975E-01 .132412991E-04    3
-.572872769E-07 .289763707E-10 .477858391E+04 .276990274E+02                   4
CYC6H9                  C   6H   9          G    300.00   5000.00 1381.00      1
 .166730638E+02 .227088190E-01-.801509353E-05 .127088484E-08-.748275111E-13    2
 .698387216E+04-.723601536E+02-.631908086E+01 .726795534E-01-.484456826E-04    3
 .157628084E-07-.202092558E-11 .153574632E+05 .524769640E+02                   4
RALDEST                 C   6H   9O   3     G    300.00   5000.00 1373.00      1
 .215153215E+02 .236419666E-01-.830694270E-05 .131026314E-08-.767602984E-13    2
-.530993462E+05-.770487448E+02 .687062608E+01 .492844450E-01-.217786396E-04    3
 .243527207E-08 .464021620E-12-.470662293E+05 .479532953E+01                   4
CYC6H11                 C   6H  11          G    300.00   5000.00 1674.00      1
 .146799252E+02 .309324453E-01-.112934485E-04 .183887582E-08-.110464203E-12    2
-.197594614E+03-.590168221E+02-.757310296E+01 .766896480E-01-.424441426E-04    3
 .941423236E-08-.439999709E-12 .764576045E+04 .620172120E+02                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   5000.00 1375.00      1
 .243899542E+02 .262326944E-01-.930434909E-05 .148019558E-08-.873538395E-13    2
-.163135893E+05-.107549099E+03-.378907832E+01 .841562901E-01-.510965662E-04    3
 .133666762E-07-.102528616E-11-.580881865E+04 .464783226E+02                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   5000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   5000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-OO                 C   6H  11O   2     G    300.00   5000.00 1380.00      1
 .225527144E+02 .280656231E-01-.990087442E-05 .156942170E-08-.923867180E-13    2
-.209455781E+05-.994788807E+02-.594021024E+01 .887171975E-01-.569424328E-04    3
 .171601250E-07-.191055830E-11-.104841379E+05 .556048484E+02                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   5000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128893429E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .565320100E+02                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   5000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   5000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
RDIPE                   C   6H  13O   1     G    300.00   5000.00 1389.00      1
 .195346832E+02 .300586517E-01-.103564671E-04 .161544621E-08-.940217507E-13    2
-.289625035E+05-.700231442E+02-.545711430E-01 .748436725E-01-.509801332E-04    3
 .191769721E-07-.313046382E-11-.218696353E+05 .358513387E+02                   4
C7H7                    C   7H   7          G    300.00   5000.00 1000.00      1
 .126890424E+02 .248754040E-01-.820402330E-05 .901804910E-09 .000000000E+00    2
 .179417186E+05-.454264236E+02-.296228400E+01 .659171040E-01-.433334430E-04    3
 .106408510E-07 .000000000E+00 .223472400E+05 .359657700E+02                   4
C6H4CH3                 C   7H   7          G    300.00   5000.00 1000.00      1
 .989521100E+01 .281997140E-01-.985390310E-05 .114532240E-08 .000000000E+00    2
 .307512908E+05-.257557742E+02-.298827000E+01 .621039310E-01-.390118950E-04    3
 .928257830E-08 .000000000E+00 .343676800E+05 .412025200E+02                   4
RCRESOLC                C   7H   7O   1     G    300.00   5000.00 1000.00      1
 .689970000E+01 .376640500E-01-.142499000E-04 .245139600E-08-.159215300E-12    2
-.104378100E+04-.796692700E+01-.415304900E+01 .776998800E-01-.583028700E-04    3
 .178677900E-07-.536299700E-12 .896696700E+03 .453288900E+02                   4
RCRESOLO                C   7H   7O   1     G    300.00   5000.00 1000.00      1
 .632623400E+01 .370920700E-01-.137369600E-04 .232847100E-08-.149701800E-12    2
-.156635900E+04-.468621100E+01-.403964400E+01 .739909500E-01-.515945300E-04    3
 .120372800E-07 .143210200E-11 .225707600E+03 .453169300E+02                   4
NC7H13                  C   7H  13          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
RMCYC6                  C   7H  13          G    300.00   5000.00 2030.00      1
 .173202469E+02 .361144629E-01-.130438584E-04 .210911191E-08-.126098895E-12    2
-.514813032E+04-.717714814E+02-.853970231E+01 .919151844E-01-.546389770E-04    3
 .144889205E-07-.127842414E-11 .374687760E+04 .679730355E+02                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   5000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
NC7H13O2                C   7H  13O   2     G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   5000.00 1386.00      1
 .252650839E+02 .325458915E-01-.113494502E-04 .178540172E-08-.104551384E-12    2
-.262255150E+05-.112686720E+03-.606776148E+01 .998265984E-01-.637962761E-04    3
 .191011484E-07-.207496071E-11-.148337709E+05 .575547331E+02                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   5000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   5000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   5000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
NC7H15                  C   7H  15          G    300.00   5000.00 1382.00      1
 .216371448E+02 .323324804E-01-.109273807E-04 .168357060E-08-.971774091E-13    2
-.105877217E+05-.852228493E+02-.379155767E-01 .756726570E-01-.407473634E-04    3
 .932678943E-08-.492360745E-12-.235605303E+04 .337321506E+02                   4
NC7H15-OO               C   7H  15O   2     G    300.00   5000.00 1393.00      1
 .272928290E+02 .327034748E-01-.112483701E-04 .175282538E-08-.101955579E-12    2
-.235449480E+05-.109307876E+03 .137396160E+01 .925294066E-01-.644403647E-04    3
 .235223293E-07-.356678305E-11-.144154775E+05 .302419431E+02                   4
NC7-QOOH                C   7H  15O   2     G    300.00   5000.00 1000.00      1
 .449365222E+02 .384325070E-02-.181753210E-06-.116055420E-10 .168632530E-14    2
-.301866739E+05-.207157897E+03 .169959950E+01 .943723540E-01-.755904260E-04    3
 .401131540E-07-.120065810E-10-.147076150E+05 .283145640E+02                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   5000.00 1395.00      1
 .269436049E+02 .351661203E-01-.120111248E-04 .186268617E-08-.107974911E-12    2
-.478858130E+05-.104588181E+03 .234060326E+01 .923428863E-01-.637138459E-04    3
 .236026902E-07-.368902757E-11-.392112217E+05 .278171493E+02                   4
C6H4C2H                 C   8H   5          G    300.00   5000.00 1000.00      1
 .286860656E+02-.138698600E-01 .227211900E-04-.998822700E-08 .140859000E-11    2
 .560473490E+05-.127502636E+03-.293242200E+01 .660436800E-01-.395005000E-04    3
-.318303810E-08 .853003870E-11 .653240430E+05 .380586850E+02                   4
C6H5C2H2                C   8H   7          G    300.00   5000.00 1394.00      1
 .187667289E+02 .200619262E-01-.690883699E-05 .107799789E-08-.627759176E-13    2
 .376789029E+05-.760287256E+02-.272251268E+01 .709701368E-01-.527526320E-04    3
 .197369835E-07-.295890798E-11 .450007235E+05 .390143531E+02                   4
RXYLENE                 C   8H   9          G    300.00   5000.00 1000.00      1
 .808697123E+01 .442230490E-01-.196920930E-04 .391313300E-08-.286780230E-12    2
 .152828351E+05-.180507988E+02-.244083000E+01 .750206000E-01-.520941000E-04    3
 .184357000E-07-.267709000E-11 .180599500E+05 .358328500E+02                   4
C8H9                    C   8H   9          G    300.00   5000.00 1000.00      1
 .179749910E+02 .239625180E-01-.715492520E-05 .103757720E-08-.596944840E-13    2
 .194242850E+05-.693345570E+02-.526520200E+01 .889877600E-01-.754492360E-04    3
 .341497320E-07-.666954430E-11 .259605610E+05 .509400020E+02                   4
RUME7                   C   8H  13O   2     G    300.00   5000.00 1376.00      1
 .270534591E+02 .305004468E-01-.106520501E-04 .167796515E-08-.983020287E-13    2
-.363346010E+05-.107800076E+03 .366021323E+01 .765652941E-01-.421034444E-04    3
 .990005395E-08-.618141131E-12-.272971814E+05 .209764369E+02                   4
RME7                    C   8H  15O   2     G    300.00   5000.00 1382.00      1
 .283088733E+02 .346001847E-01-.117889297E-04 .182346779E-08-.105527368E-12    2
-.507031223E+05-.115791454E+03 .312712425E+01 .886538094E-01-.550709022E-04    3
 .172495936E-07-.218153163E-11-.414147165E+05 .212562509E+02                   4
IC8H17                  C   8H  17          G    300.00   5000.00 1000.00      1
 .210071027E+02 .400670210E-01-.122220840E-04 .179139180E-08-.103364050E-12    2
-.156827594E+05-.841376688E+02-.142527150E+01 .952433870E-01-.515412500E-04    3
 .269038680E-08 .557281520E-11-.909216410E+04 .335841900E+02                   4
IC8H17-OO               C   8H  17O   2     G    300.00   5000.00 1397.00      1
 .307492955E+02 .368544999E-01-.126522533E-04 .196915974E-08-.114442369E-12    2
-.380116818E+05-.129042218E+03-.126574300E+01 .113828908E+00-.844050615E-04    3
 .328104935E-07-.525271208E-11-.270886887E+05 .421608430E+02                   4
IC8-QOOH                C   8H  17O   2     G    300.00   5000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   5000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   5000.00 1398.00      1
 .362956073E+02 .372755603E-01-.128091685E-04 .199516372E-08-.116026947E-12    2
-.507708950E+05-.153592254E+03 .134208862E+01 .119507370E+00-.864939904E-04    3
 .319097725E-07-.475802942E-11-.387629197E+05 .338018650E+02                   4
INDENYL                 C   9H   7          G    300.00   5000.00 1389.00      1
 .210619876E+02 .219045968E-01-.772700080E-05 .122481766E-08-.721012249E-13    2
 .270100509E+05-.947705468E+02-.627808779E+01 .881610767E-01-.698280991E-04    3
 .280009421E-07-.454051640E-11 .362473103E+05 .511874555E+02                   4
RC9H11                  C   9H  11          G    300.00   5000.00 1385.00      1
 .227307929E+02 .291439937E-01-.101635526E-04 .159859987E-08-.935933623E-13    2
 .481056390E+04-.975266902E+02-.180604559E+01 .826070356E-01-.539943357E-04    3
 .177716542E-07-.237645289E-11 .137819561E+05 .357292291E+02                   4
C10H7                   C  10H   7          G    300.00   5000.00 1000.00      1
 .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
 .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
 .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
C10H7O                  C  10H   7O   1     G    300.00   5000.00 1387.00      1
 .252263199E+02 .234793777E-01-.827533154E-05 .131107385E-08-.771548491E-13    2
 .188945294E+04-.112699321E+03-.234081413E+01 .850055448E-01-.590412510E-04    3
 .195981954E-07-.248272174E-11 .116463286E+05 .362009562E+02                   4
RTETRALIN               C  10H  11          G    300.00   5000.00 1393.00      1
 .274897602E+02 .290231662E-01-.101643070E-04 .160474752E-08-.942455736E-13    2
 .498834588E+04-.134140516E+03-.103201226E+02 .112759920E+00-.777366610E-04    3
 .248527119E-07-.289510552E-11 .183518811E+05 .701782401E+02                   4
RTETRAOO                C  10H  11O   2     G    300.00   5000.00 1393.00      1
 .325696052E+02 .270322587E-01-.103226960E-04 .172977036E-08-.105947326E-12    2
-.797598133E+04-.153101057E+03-.133437809E+02 .139730780E+00-.110918062E-03    3
 .406822937E-07-.565600132E-11 .639529388E+04 .899902305E+02                   4
RDECALIN                C  10H  17          G    300.00   5000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
RODECA                  C  10H  17          G    300.00   5000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
QDECOOH                 C  10H  17O   2     G    300.00   5000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
RDECOO                  C  10H  17O   2     G    300.00   5000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
ZDECA                   C  10H  17O   4     G    300.00   5000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
NC10H19                 C  10H  19          G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC10H19O2               C  10H  19O   2     G    300.00   5000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC10H21                 C  10H  21          G    300.00   5000.00 1385.00      1
 .314447580E+02 .452778532E-01-.153145696E-04 .236072411E-08-.136311835E-12    2
-.229702700E+05-.131435127E+03-.930536886E+00 .113137924E+00-.664034118E-04    3
 .183220872E-07-.177128003E-11-.109890165E+05 .451328034E+02                   4
NC10-QOOH               C  10H  21O   2     G    300.00   5000.00 1392.00      1
 .364873664E+02 .456938220E-01-.154604572E-04 .238346695E-08-.137626430E-12    2
-.370093465E+05-.152798812E+03 .883511244E+00 .125360621E+00-.820308363E-04    3
 .270294818E-07-.354081617E-11-.243570772E+05 .395546233E+02                   4
NC10H21-OO              C  10H  21O   2     G    300.00   5000.00 1392.00      1
 .347424373E+02 .481682266E-01-.165183738E-04 .256870455E-08-.149189141E-12    2
-.416206773E+05-.145293449E+03 .109633829E+01 .123998092E+00-.822926235E-04    3
 .288935474E-07-.426829326E-11-.295195291E+05 .366210584E+02                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   5000.00 1393.00      1
 .419701067E+02 .470326141E-01-.162065055E-04 .252885796E-08-.147242779E-12    2
-.568721943E+05-.179987435E+03 .270340236E+01 .134161981E+00-.884509572E-04    3
 .291143638E-07-.380678318E-11-.428023111E+05 .324857210E+02                   4
C10H6CH3                C  11H   9          G    300.00   5000.00 1387.00      1
 .241866524E+02 .287085863E-01-.100040198E-04 .157283341E-08-.920615442E-13    2
 .317595121E+05-.107209439E+03-.148986180E+01 .837301572E-01-.531437515E-04    3
 .161159556E-07-.183550466E-11 .411521411E+05 .324161445E+02                   4
C10H7CH2                C  11H   9          G    300.00   5000.00 1389.00      1
 .266596927E+02 .269903845E-01-.949827903E-05 .150313533E-08-.883831941E-13    2
 .210179470E+05-.122975754E+03-.551514480E+01 .106245066E+00-.857510752E-04    3
 .355122444E-07-.598055713E-11 .318146452E+05 .484291679E+02                   4
CH3C10H6O               C  11H   9O   1     G    300.00   5000.00 1386.00      1
 .281108749E+02 .281427040E-01-.986090177E-05 .155620703E-08-.913337710E-13    2
-.350666986E+04-.125748079E+03-.108570461E+01 .905308669E-01-.577474885E-04    3
 .167977934E-07-.168045736E-11 .709977655E+04 .329292729E+02                   4
RUME10                  C  11H  19O   2     G    300.00   5000.00 1400.00      1
 .333201898E+02 .479399831E-01-.157699228E-04 .238393079E-08-.135735725E-12    2
-.400970534E+05-.137405141E+03 .142231026E+01 .127120401E+00-.922642215E-04    3
 .364453822E-07-.599028369E-11-.294852312E+05 .322500169E+02                   4
RMDX                    C  11H  21O   2     G    300.00   5000.00 1376.00      1
 .385051195E+02 .464902832E-01-.162008540E-04 .254969816E-08-.149299808E-12    2
-.649901621E+05-.166525707E+03 .345128941E+01 .114960511E+00-.621890037E-04    3
 .140937438E-07-.752795690E-12-.513892174E+05 .266431624E+02                   4
RMDOOX                  C  11H  21O   4     G    300.00   5000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
QMDOOH                  C  11H  21O   4     G    300.00   5000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
ZMDOOH                  C  11H  21O   6     G    300.00   5000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
C12H7                   C  12H   7          G    300.00   5000.00 1000.00      1
 .119534365E+02 .523860720E-01-.276952580E-04 .698583900E-08-.684938540E-12    2
 .531995141E+05-.403925438E+02-.733802700E+01 .111965800E+00-.932829430E-04    3
 .358663430E-07-.426602200E-11 .580597660E+05 .573507160E+02                   4
RBIPHENYL               C  12H   9          G    300.00   5000.00 1000.00      1
 .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
 .415521488E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
 .194042280E-07 .000000000E+00 .498170300E+05 .608493300E+02                   4
NC12H25                 C  12H  25          G    300.00   5000.00 1387.00      1
 .379559371E+02 .541231481E-01-.184408520E-04 .285618139E-08-.165452331E-12    2
-.312698454E+05-.166157365E+03-.117025753E+01 .136564242E+00-.813840519E-04    3
 .231564976E-07-.240764498E-11-.167979250E+05 .471339366E+02                   4
NC12-QOOH               C  12H  25O   2     G    300.00   5000.00 1392.00      1
 .427882927E+02 .547351985E-01-.185693137E-04 .286771608E-08-.165782124E-12    2
-.451897912E+05-.183774591E+03 .457142729E+00 .149660990E+00-.984019129E-04    3
 .327982507E-07-.438634589E-11-.301386488E+05 .448987214E+02                   4
NC12H25-OO              C  12H  25O   2     G    300.00   5000.00 1392.00      1
 .410672882E+02 .571682582E-01-.196096581E-04 .304996352E-08-.177163659E-12    2
-.498119415E+05-.176403781E+03 .761653139E+00 .147870053E+00-.980093227E-04    3
 .342486611E-07-.502171364E-11-.353144020E+05 .415448990E+02                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   5000.00 1393.00      1
 .478223133E+02 .563342752E-01-.193784199E-04 .302016363E-08-.175696376E-12    2
-.648031378E+05-.208209874E+03 .250560092E+01 .157994999E+00-.105503812E-03    3
 .358709948E-07-.494871123E-11-.486270464E+05 .366890378E+02                   4
C14H9                   C  14H   9          G    300.00   5000.00 1000.00      1
 .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
 .431324738E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
 .240156710E-07 .000000000E+00 .527750200E+05 .639753600E+02                   4
C16H9                   C  16H   9          G    300.00   5000.00 1000.00      1
 .161628784E+02 .696969850E-01-.371786410E-04 .946306230E-08-.935417110E-12    2
 .461067047E+05-.652717249E+02-.114972670E+02 .151166960E+00-.116351410E-03    3
 .317097570E-07 .218082760E-11 .532378630E+05 .757195740E+02                   4
IC16H33                 C  16H  33          G    300.00   5000.00 1398.00      1
 .560389730E+02 .668182464E-01-.225681513E-04 .347608102E-08-.200620637E-12    2
-.583645424E+05-.270643351E+03-.953227198E+01 .224283987E+00-.166371012E-03    3
 .627848165E-07-.951119300E-11-.362947496E+05 .795385858E+02                   4
NC16H33                 C  16H  33          G    300.00   5000.00 1387.00      1
 .510324990E+02 .711045684E-01-.240491592E-04 .370710805E-08-.214054039E-12    2
-.477151440E+05-.228063103E+03-.243005348E+01 .186692969E+00-.115724867E-03    3
 .350879669E-07-.405848895E-11-.282942913E+05 .622394761E+02                   4
IC16H33-OO              C  16H  33O   2     G    300.00   5000.00 1397.00      1
 .600009189E+02 .697612153E-01-.240119992E-04 .374399505E-08-.217877031E-12    2
-.771125672E+05-.288496873E+03-.807177622E+01 .238256241E+00-.186291159E-03    3
 .758296536E-07-.125956694E-10-.544214916E+05 .737310481E+02                   4
NC16H33-OO              C  16H  33O   2     G    300.00   5000.00 1392.00      1
 .537254976E+02 .751675700E-01-.257930312E-04 .401271756E-08-.233130903E-12    2
-.661992854E+05-.238675214E+03 .121036107E+00 .195526928E+00-.129332034E-03    3
 .448994551E-07-.651714304E-11-.469097176E+05 .512502917E+02                   4
NC16-QOOH               C  16H  33O   2     G    300.00   5000.00 1394.00      1
 .557196631E+02 .758805933E-01-.260092776E-04 .404350192E-08-.234807139E-12    2
-.852319237E+05-.250905152E+03-.858601178E+00 .204663464E+00-.138309577E-03    3
 .488963438E-07-.717831502E-11-.651200924E+05 .543621098E+02                   4
IC16-QOOH               C  16H  33O   2     G    300.00   5000.00 1399.00      1
 .615798034E+02 .683372119E-01-.235040286E-04 .366308625E-08-.213104512E-12    2
-.710887760E+05-.294961987E+03-.836284759E+01 .243137667E+00-.193204766E-03    3
 .794478202E-07-.132585716E-10-.480052296E+05 .765156723E+02                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   5000.00 1397.00      1
 .619590914E+02 .670805941E-01-.228781110E-04 .354645272E-08-.205581639E-12    2
-.737750910E+05-.297686975E+03-.828638110E+01 .240615134E+00-.188046280E-03    3
 .753924180E-07-.122092604E-10-.505105835E+05 .759168895E+02                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   5000.00 1393.00      1
 .605564321E+02 .743085731E-01-.255622121E-04 .398394439E-08-.231762903E-12    2
-.812450313E+05-.270973587E+03 .185761468E+01 .205470409E+00-.136236709E-03    3
 .460471713E-07-.632675050E-11-.602164277E+05 .464682670E+02                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   5000.00 1396.00      1
 .664600695E+02 .692200495E-01-.239811044E-04 .375550159E-08-.219211037E-12    2
-.927495777E+05-.318609160E+03-.734744585E+01 .256652224E+00-.210530384E-03    3
 .896944245E-07-.155165690E-10-.685533247E+05 .725686554E+02                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   5000.00 1395.00      1
 .657312368E+02 .698159219E-01-.241818212E-04 .378635278E-08-.220988765E-12    2
-.891725518E+05-.313140345E+03-.709314164E+01 .252307521E+00-.202956898E-03    3
 .848048060E-07-.144255682E-10-.650715559E+05 .736645741E+02                   4
RUME16                  C  17H  31O   2     G    300.00   5000.00 1836.00      1
 .492312959E+02 .809629787E-01-.290414743E-04 .466984560E-08-.277987170E-12    2
-.712766099E+05-.212350222E+03 .581847898E+00 .197335153E+00-.132222747E-03    3
 .454132116E-07-.638160297E-11-.555076491E+05 .468001664E+02                   4
RMPAX                   C  17H  33O   2     G    300.00   5000.00 1000.00      1
 .347969412E+02 .108174887E+00-.436560662E-04 .805036686E-08-.557001848E-12    2
-.833532968E+05-.136711346E+03 .118429649E+02 .108281798E+00 .937470576E-04    3
-.175260710E-06 .681980157E-10-.741770519E+05-.304443036E+01                   4
QMPAOOH                 C  17H  33O   4     G    300.00   5000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
RMPAOOX                 C  17H  33O   4     G    300.00   5000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   5000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
RMLIN1X                 C  19H  31O   2     G    300.00   5000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1A                 C  19H  31O   2     G    300.00   5000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   5000.00 1854.00      1
 .566771062E+02 .848718923E-01-.306165992E-04 .494186779E-08-.294961213E-12    2
-.712260452E+05-.243221478E+03-.182318626E+01 .229267759E+00-.163619600E-03    3
 .597071790E-07-.884702825E-11-.526983896E+05 .668009912E+02                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   5000.00 1859.00      1
 .597198037E+02 .825172318E-01-.298594827E-04 .482987333E-08-.288709215E-12    2
-.679692648E+05-.260058551E+03-.300959205E+01 .239625356E+00-.176824958E-03    3
 .662378545E-07-.999748235E-11-.483423909E+05 .715224170E+02                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   5000.00 1844.00      1
 .633953698E+02 .840133680E-01-.304696355E-04 .493592631E-08-.295352525E-12    2
-.861431583E+05-.275575442E+03 .377427203E+00 .239045319E+00-.172299424E-03    3
 .627369839E-07-.920510825E-11-.661691485E+05 .585014961E+02                   4
RMLINX                  C  19H  33O   2     G    300.00   5000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLINA                  C  19H  33O   2     G    300.00   5000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLINOOX                C  19H  33O   4     G    300.00   5000.00 1840.00      1
 .561396497E+02 .898573320E-01-.323076347E-04 .520295879E-08-.310043109E-12    2
-.835647272E+05-.240835194E+03 .146002415E+01 .221120424E+00-.149309126E-03    3
 .517229930E-07-.733489301E-11-.658774535E+05 .502873652E+02                   4
QMLINOOX                C  19H  33O   4     G    300.00   5000.00 1830.00      1
 .592334771E+02 .871071695E-01-.313329462E-04 .504827960E-08-.300945381E-12    2
-.780101129E+05-.256778117E+03-.383425349E+00 .231626065E+00-.160960610E-03    3
 .566395921E-07-.805109149E-11-.589322117E+05 .599912602E+02                   4
ZMLINOOX                C  19H  33O   6     G    300.00   5000.00 1183.00      1
 .601829822E+02 .877246704E-01-.308673874E-04 .490011538E-08-.289106438E-12    2
-.959756017E+05-.274111539E+03 .888177201E+00 .245491279E+00-.188867182E-03    3
 .756398491E-07-.122061299E-10-.781464330E+05 .361650421E+02                   4
RMEOLES                 C  19H  35O   2     G    300.00   5000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLEA                 C  19H  35O   2     G    300.00   5000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   5000.00 1799.00      1
 .565118676E+02 .949710722E-01-.342666750E-04 .553134168E-08-.330143553E-12    2
-.121723087E+06-.240377715E+03 .312228984E+01 .215930145E+00-.133878272E-03    3
 .413627115E-07-.514696341E-11-.103763030E+06 .464356398E+02                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   5000.00 1000.00      1
 .578903822E+02 .960618008E-01-.345783142E-04 .557312937E-08-.332293982E-12    2
-.145787244E+06-.248797880E+03-.121085721E+01 .236084007E+00-.157011163E-03    3
 .530523572E-07-.729693062E-11-.126516243E+06 .664772594E+02                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   5000.00 1000.00      1
 .558298346E+02 .101939581E+00-.350749088E-04 .548251413E-08-.319925836E-12    2
-.108843753E+06-.228788516E+03 .196924109E+01 .244903891E+00-.177892306E-03    3
 .692918136E-07-.110530115E-10-.926192007E+05 .531689573E+02                   4
RSTEAX                  C  19H  37O   2     G    300.00   5000.00 1000.00      1
 .410838828E+02 .116388491E+00-.460844475E-04 .839784976E-08-.576703150E-12    2
-.912925804E+05-.167019971E+03 .115570681E+02 .131479341E+00 .799583356E-04    3
-.171755777E-06 .679701047E-10-.799964069E+05 .174630364E+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   5000.00 1384.00      1
 .294145201E+02 .809900030E-01-.261520592E-04 .393935978E-08-.226643615E-12    2
-.317656348E+05-.119394359E+03 .329283081E+01 .226000653E+00-.143515509E-03    3
 .442428385E-07-.517811632E-11-.232845416E+05 .214592368E+02                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   5000.00 1378.00      1
 .297828900E+02 .771449164E-01-.253926493E-04 .388430700E-08-.225914471E-12    2
-.317651562E+05-.119207488E+03 .391542481E+01 .223377046E+00-.136351584E-03    3
 .377005603E-07-.345802861E-11-.232839019E+05 .214376580E+02                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   5000.00 1384.00      1
 .300794787E+02 .502955745E-01-.168090526E-04 .259970193E-08-.151164888E-12    2
-.397961494E+04-.130229963E+02 .598820430E+01 .157430576E+00-.110701951E-03    3
 .400055584E-07-.590540707E-11-.291813417E+04 .432758910E+01                   4
AC3H4                   C   3H   4          G    300.00   3500.00 1800.00      1
 6.64430238e+00 1.14987825e-02-4.68099585e-06 9.62334222e-10-8.24360065e-14    2
 2.07131189e+04-1.35744541e+01 1.21562918e+00 2.35625008e-02-1.47340944e-05    3
 4.68570404e-09-5.99570704e-13 2.26674413e+04 1.58066578e+01                   4
ACETOL                  C   3H   6O   2     G    300.00   3500.00 1800.00      1
 9.43106557e+00 1.86879303e-02-7.29283976e-06 1.39932581e-09-1.08736168e-13    2
-4.87389994e+04-2.08360480e+01 1.41553145e+00 3.65002283e-02-2.21364215e-05    3
 6.89694866e-09-8.72294898e-13-4.58534071e+04 2.25456947e+01                   4
ALDEST                  C   6H  10O   3     G    300.00   3500.00 1800.00      1
 1.79608805e+01 3.27577303e-02-1.29904809e-05 2.50013680e-09-1.93431386e-13    2
-7.48983193e+04-5.99171462e+01 5.24137808e+00 6.10232913e-02-3.65451150e-05    3
 1.12240754e-08-1.40508952e-12-7.03192984e+04 8.92345431e+00                   4
ALDINS                  C  13H  20O   1     G    300.00   3500.00 1800.00      1
 8.44295858e+01 4.93170400e-02-2.86268350e-05 8.86979917e-09-1.00373619e-12    2
-8.94265291e+04-4.12065762e+02-1.18024916e+01 2.63166101e-01-2.06834386e-04    3
 7.48725957e-08-1.01707913e-11-5.47829813e+04 1.08762316e+02                   4
AR                      AR  1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
-7.45375000e+02 4.36600000e+00 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25-7.45375000e+02 4.36600000e+00                   4
BENZYNE                 C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465819e+01 1.50373246e-02-5.27844959e-06 8.14607581e-10-4.49073366e-14    2
 5.03301418e+04-3.53782934e+01-3.73796173e+00 5.69931634e-02-5.02311341e-05    3
 2.22206478e-08-3.86741452e-12 5.44418140e+04 4.04070822e+01                   4
BIN1A                   C  20H  16          G    300.00   3500.00 1800.00      1
-3.24173600e+00 1.58222900e-01-9.46183500e-05 2.81843100e-08-3.56131000e-12    2
 2.17869900e+04 3.00825300e+01-3.24173600e+00 1.58222900e-01-9.46183500e-05    3
 2.81843100e-08-3.56131000e-12 2.17869900e+04 3.00825300e+01                   4
BIN1B                   C  20H  10          G    300.00   3500.00 1800.00      1
-5.70256700e+00 1.43432300e-01-8.80724700e-05 2.76799200e-08-3.52289900e-12    2
 2.77808900e+04 4.34481200e+01-5.70256700e+00 1.43432300e-01-8.80724700e-05    3
 2.76799200e-08-3.52289900e-12 2.77808900e+04 4.34481200e+01                   4
BIPHENYL                C  12H  10          G    300.00   3500.00 1450.00      1
 2.67692078e+01 2.81611415e-02-6.05667723e-06-3.69378426e-10 1.67249382e-13    2
 9.26692468e+03-1.21306413e+02-1.05625108e+01 1.31145193e-01-1.12591903e-04    3
 4.86123345e-08-8.27787353e-12 2.00931231e+04 7.26686556e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623567e-02-8.52218599e-06 1.36123710e-09-7.97159891e-14    2
-5.90596972e+03-6.59480381e+01-8.70136947e+00 9.66875823e-02-8.77887356e-05    3
 3.96542562e-08-7.01685714e-12 1.03797027e+03 6.35339364e+01                   4
C                       C   1               G    300.00   3500.00  700.00      1
 2.48989675e+00 5.14965671e-05-7.37912415e-08 3.75721674e-11-4.86583734e-15    2
 8.54527782e+04 4.81783270e+00 2.55088394e+00-2.97001640e-04 6.72990632e-07    3
-6.73648664e-10 2.49141603e-13 8.54442400e+04 4.54535738e+00                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934216e-02-1.83631832e-05 3.88491136e-09-3.27420808e-13    2
 4.39687821e+03-8.23923218e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836942e-12 1.50954180e+04 7.84485932e+01                   4
C10H6CH3                C  11H   9          G    300.00   3500.00 1800.00      1
 2.12659882e+01 3.44429430e-02-1.39605695e-05 2.72496148e-09-2.12674976e-13    2
 3.28507521e+04-9.11529083e+01-1.92673037e+00 8.59823175e-02-5.69100482e-05    3
 1.86321758e-08-2.42201030e-12 4.12001308e+04 3.43709226e+01                   4
C10H7                   C  10H   7          G    300.00   3500.00 1440.00      1
 1.86034915e+01 2.84557463e-02-7.51492092e-06 8.59843958e-11 1.31843536e-13    2
 3.89175328e+04-7.96671600e+01-8.11601745e+00 1.02676605e-01-8.48283149e-05    3
 3.58792224e-08-6.08226028e-12 4.66127513e+04 5.89821104e+01                   4
C10H7CH2                C  11H   9          G    300.00   3500.00 1460.00      1
 1.62958766e+01 4.54296741e-02-2.13529357e-05 4.77934912e-09-4.18010504e-13    2
 2.55100815e+04-6.47739136e+01-5.20583638e+00 1.04338477e-01-8.18756782e-05    3
 3.24153046e-08-5.15019466e-12 3.17885817e+04 4.70964540e+01                   4
C10H7CH3                C  11H  10          G    300.00   3500.00 1400.00      1
 1.59718633e+01 4.84656090e-02-2.27123224e-05 5.09437338e-09-4.47432797e-13    2
 5.32412011e+03-6.35417268e+01-7.85505905e+00 1.16542530e-01-9.56518805e-05    3
 3.98274963e-08-6.64977617e-12 1.19956584e+04 5.94264980e+01                   4
C10H7CHO                C  11H   8O   1     G    300.00   3500.00 1800.00      1
 2.76873866e+01 2.65153545e-02-9.85230690e-06 1.73492056e-09-1.21699947e-13    2
-1.08926269e+04-1.25645702e+02-1.80645208e+00 9.20572182e-02-6.44705267e-05    3
 2.19638908e-08-2.93127915e-12-2.74844971e+02 3.39811053e+01                   4
C10H7O                  C  10H   7O   1     G    300.00   3500.00 1800.00      1
 2.60845785e+01 2.24488808e-02-7.86244785e-06 1.25147148e-09-7.55452008e-14    2
 1.36168392e+03-1.17834769e+02-2.53985295e+00 8.60587284e-02-6.08706542e-05    3
 2.08841405e-08-2.80230479e-12 1.16664792e+04 3.70866255e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248659e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987876e+01                   4
C11H12O4                C  11H  12O   4     G    300.00   3500.00 1280.00      1
 2.98957517e+01 4.73870505e-02-2.11603212e-05 4.60350399e-09-3.96349099e-13    2
-7.02119467e+04-1.21160681e+02-3.09348688e+00 1.50478421e-01-1.41970521e-04    3
 6.75254832e-08-1.26857982e-11-6.17667016e+04 4.61370519e+01                   4
C12H18                  C  12H  18          G    300.00   3500.00 1800.00      1
 8.44295858e+01 4.93170400e-02-2.86268350e-05 8.86979917e-09-1.00373619e-12    2
-8.94265291e+04-4.12065762e+02-1.18024916e+01 2.63166101e-01-2.06834386e-04    3
 7.48725957e-08-1.01707913e-11-5.47829813e+04 1.08762316e+02                   4
C12H22                  C  12H  22          G    300.00   3500.00 1760.00      1
 3.60687856e+01 4.93531801e-02-1.68932777e-05 2.64866878e-09-1.56934744e-13    2
-2.29291143e+04-1.58689972e+02-2.71855262e+00 1.37506222e-01-9.20237107e-05    3
 3.11071661e-08-4.19933494e-12-9.27597128e+03 5.03635315e+01                   4
C12H7                   C  12H   7          G    300.00   3500.00 1250.00      1
 1.23349807e+01 5.16907682e-02-2.72404819e-05 6.85858162e-09-6.72018930e-13    2
 5.30394981e+04-4.25244963e+01-8.02968441e+00 1.16857696e-01-1.05440796e-04    3
 4.85654157e-08-9.01338574e-12 5.81306643e+04 6.02674845e+01                   4
C12H8                   C  12H   8          G    300.00   3500.00 1430.00      1
 2.59652189e+01 2.42501190e-02-4.81412894e-06-4.21078741e-10 1.47447105e-13    2
 1.90778575e+04-1.18254954e+02-9.28199067e+00 1.22843712e-01-1.08233982e-04    3
 4.77933050e-08-8.28164096e-12 2.91585594e+04 6.43994840e+01                   4
C14H10                  C  14H  10          G    300.00   3500.00 1430.00      1
 3.13141255e+01 2.89528714e-02-5.57670990e-06-5.89662906e-10 1.88202945e-13    2
 1.06460191e+04-1.48101025e+02-1.21905872e+01 1.50644375e-01-1.33225141e-04    3
 5.89200950e-08-1.02156009e-11 2.30883669e+04 7.73445897e+01                   4
C14H9                   C  14H   9          G    300.00   3500.00 1430.00      1
 3.13141255e+01 2.89528714e-02-5.57670990e-06-5.89662906e-10 1.88202945e-13    2
 4.06560892e+04-1.48101025e+02-1.21905872e+01 1.50644375e-01-1.33225141e-04    3
 5.89200950e-08-1.02156009e-11 5.30984370e+04 7.73445897e+01                   4
C16H10                  C  16H  10          G    300.00   3500.00 1430.00      1
 3.55205969e+01 2.97059226e-02-5.18577408e-06-7.74976601e-10 2.05764301e-13    2
 1.13998034e+04-1.72584653e+02-1.43149515e+01 1.69106058e-01-1.51409692e-04    3
 6.73946823e-08-1.17120082e-11 2.56527702e+04 8.56679628e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933977e+01 6.96117135e-02-3.71054121e-05 9.43826014e-09-9.32515880e-13    2
 4.61008358e+04-6.54256237e+01-1.33382684e+01 1.64875153e-01-1.52343443e-04    3
 7.13941909e-08-1.34236310e-11 5.34246890e+04 8.34001920e+01                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319129e-02-1.90892866e-05    3
 5.92848300e-09-7.42884555e-13-1.63833552e+04 6.70139036e+00                   4
C2-OQOOH                C   2H   4O   3     G    300.00   3500.00 1800.00      1
 1.06961666e+01 1.25934013e-02-5.32391821e-06 1.08565058e-09-8.80671200e-14    2
-3.42000230e+04-2.43964294e+01 5.53941294e+00 2.40528540e-02-1.48734621e-05    3
 4.62251869e-09-5.79298801e-13-3.23435917e+04 3.51299738e+00                   4
C2-QOOH                 C   2H   5O   2     G    300.00   3500.00 1270.00      1
 7.85685775e+00 1.67911217e-02-7.79621720e-06 1.73782470e-09-1.51982948e-13    2
 7.20248835e+02-1.06887184e+01 8.24295798e-01 3.89409231e-02-3.39574000e-05    3
 1.54707291e-08-2.85531058e-12 2.50651957e+03 2.49202290e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1770.00      1
 2.62706056e+00 5.61439161e-03-2.33738366e-06 4.29433761e-10-2.92352464e-14    2
 6.73836200e+04 9.73315238e+00 4.71151838e+00 9.03752455e-04 1.65468342e-06    3
-1.07416966e-09 1.83138118e-13 6.66457220e+04-1.51333448e+00                   4
C2H2                    C   2H   2          G    300.00   3500.00  970.00      1
 4.61193612e+00 5.01498204e-03-1.65253694e-06 2.49922532e-10-1.30568636e-14    2
 2.56043843e+04-3.75517096e+00 1.83812159e+00 1.64533925e-02-1.93408005e-05    3
 1.24068047e-08-3.14627391e-12 2.61425043e+04 9.54239252e+00                   4
C2H2O2                  C   2H   2O   2     G    300.00   3500.00 1700.00      1
 9.83116579e+00 4.87360532e-03-1.69443300e-06 2.65361078e-10-1.54439841e-14    2
-2.96273239e+04-2.66407027e+01 1.89947966e+00 2.35363962e-02-1.81616014e-05    3
 6.72307419e-09-9.65107677e-13-2.69305506e+04 1.58338747e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00  700.00      1
 7.05094230e-01 1.53761148e-02-8.91788178e-06 2.51340905e-09-2.70561650e-13    2
 3.36189510e+04 1.96531878e+01 2.74606708e+00 3.71341276e-03 1.60736225e-05    3
-2.12880236e-08 8.22995002e-12 3.33332148e+04 1.05346375e+01                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1340.00      1
 6.70517760e+00 1.61222451e-02-7.57298869e-06 1.70307233e-09-1.49924851e-13    2
-1.33618589e+04-9.88613663e+00 3.40917666e-01 3.51200360e-02-2.88391725e-05    3
 1.22832633e-08-2.12384107e-12-1.16562372e+04 2.26803642e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1800.00      1
 4.49333672e+00 1.00335105e-02-3.62601388e-06 5.97613541e-10-3.65481279e-14    2
 3.93220822e+03-3.35192020e+00 2.66161697e-01 1.94272328e-02-1.14541158e-05    3
 3.49691054e-09-4.39228267e-13 5.45399123e+03 1.95264329e+01                   4
C2H4O                   C   2H   4O   1     G    300.00   3500.00 1440.00      1
 4.77217531e+00 1.29608883e-02-4.19608017e-06 3.32859470e-10 2.97428516e-14    2
-8.91054882e+03-2.99568268e+00-1.76683146e+00 3.11247960e-02-2.31168173e-05    3
 9.09246001e-09-1.49102113e-12-7.02731487e+03 3.09356489e+01                   4
C2H4O2                  C   2H   4O   2     G    300.00   3500.00  770.00      1
 3.40614010e+00 2.02613044e-02-1.03463461e-05 2.53497107e-09-2.40436915e-13    2
-3.88060356e+04 1.20569218e+01 4.64403525e+00 1.38306802e-02 2.18084389e-06    3
-8.31108086e-09 3.28100852e-12-3.89966715e+04 6.40833543e+00                   4
C2H4OH                  C   2H   5O   1     G    300.00   3500.00 1800.00      1
 6.43071837e+00 1.30529032e-02-5.04234033e-06 9.42421880e-10-7.06192378e-14    2
-6.84254175e+03-6.40643970e+00 1.19058412e+00 2.46976460e-02-1.47462926e-05    3
 4.53647829e-09-5.69793739e-13-4.95609342e+03 2.19542600e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00  700.00      1
-1.10489358e+00 2.43511913e-02-1.39613152e-05 3.89870297e-09-4.17285120e-13    2
 1.35030749e+04 3.00146907e+01 4.99501831e+00-1.05054480e-02 6.07314834e-05    3
-6.72372957e-08 2.49884287e-11 1.26490872e+04 2.76182763e+00                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1140.00      1
-3.19796156e+00 4.17401347e-02-2.22156952e-05 5.37596466e-09-4.95601240e-13    2
-2.31457657e+04 4.43385409e+01 4.65967589e+00 1.41694770e-02 1.40614860e-05    3
-1.58387612e-08 4.15675092e-12-2.49373071e+04 5.40040975e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1380.00      1
 4.82959470e+00 1.77552121e-02-6.21112100e-06 6.58265206e-10 1.60136692e-14    2
-3.08658494e+04 5.43180378e-01 2.48921589e-01 3.10325255e-02-2.06429833e-05    3
 7.63017938e-09-1.24701426e-12-2.96015836e+04 2.41176395e+01                   4
C2H5OO                  C   2H   5O   2     G    300.00   3500.00 1260.00      1
 4.82335647e+00 2.06819188e-02-9.67611879e-06 2.17589519e-09-1.91914821e-13    2
-4.75156327e+03 3.93765088e+00 1.82119985e+00 3.02125747e-02-2.10221378e-05    3
 8.17907984e-09-1.38302289e-12-3.99501980e+03 1.91151548e+01                   4
C2H5OOH                 C   2H   6O   2     G    300.00   3500.00 1590.00      1
 1.15652199e+01 1.02216474e-02-1.86630047e-06-2.55692055e-10 7.26211298e-14    2
-2.47328137e+04-3.42112965e+01 1.46294225e+00 3.56361824e-02-2.58422768e-05    3
 9.79712822e-09-1.50801099e-12-2.15202894e+04 1.92111233e+01                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.39373503e+00 1.52684734e-02-5.82725051e-06 1.10377088e-09-8.60486537e-14    2
-1.27269866e+04-3.21997495e+00-2.74461309e-01 2.56422430e-02-1.44720586e-05    3
 4.30555164e-09-5.30740425e-13-1.10464360e+04 2.20452775e+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   3500.00 1350.00      1
 1.12132537e+01 2.34709018e-02-1.13098317e-05 2.59008079e-09-2.30885268e-13    2
-3.91289882e+04-2.66260028e+01 8.46220448e-01 5.41880374e-02-4.54399824e-05    3
 1.94444762e-08-3.35206960e-12-3.63298893e+04 2.65001343e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00  700.00      1
 6.27665898e+00 5.58433105e-03-2.45857473e-06 5.41223006e-10-4.83608105e-14    2
 6.31055207e+04-4.75111128e+00 4.26055345e+00 1.71049341e-02-2.71455812e-05    3
 2.40526578e-08-8.44530180e-12 6.33877755e+04 4.25633816e+00                   4
C3H3                    C   3H   3          G    300.00   3500.00 1720.00      1
 1.09930471e+01 7.79714852e-04 1.73957383e-06-7.95864951e-10 9.69732207e-14    2
 3.74627231e+04-3.40822737e+01 3.56039712e+00 1.80649474e-02-1.33347569e-05    3
 5.04689889e-09-7.52265710e-13 4.00195547e+04 5.80687271e+00                   4
C3H4O2                  C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920429e+01 1.38871300e-02-6.12561993e-06 1.30548845e-09-1.09965765e-13    2
-3.57026988e+04-2.69350036e+01 1.17378045e-01 4.67086294e-02-4.58290467e-05    3
 2.26514168e-08-4.41358036e-12-3.31793820e+04 2.43405589e+01                   4
C3H4O3                  C   3H   4O   3     G    300.00   3500.00 1710.00      1
 1.37242810e+01 1.08811110e-02-3.70124855e-06 5.78901440e-10-3.43205818e-14    2
-5.77802807e+04-3.99570073e+01 2.17563103e+00 3.78954970e-02-2.73980784e-05    3
 9.81743159e-09-1.38498288e-12-5.38306424e+04 2.19543274e+01                   4
C3H5CHO                 C   4H   6O   1     G    300.00   3500.00 1610.00      1
 9.36564259e+00 1.99394689e-02-8.24714277e-06 1.63840913e-09-1.29181894e-13    2
-1.44293663e+04-2.07054000e+01 2.40474771e-01 4.26106933e-02-2.93694015e-05    3
 1.03846860e-08-1.48729943e-12-1.14910622e+04 2.76639767e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00  820.00      1
 2.45863176e+00 2.66446458e-02-1.24879759e-05 2.92198798e-09-2.71872686e-13    2
-1.72239991e+04 1.83830345e+01 4.24999286e+00 1.79062989e-02 3.49680492e-06    3
-1.00737688e-08 3.69024828e-12-1.75177823e+04 1.00962500e+01                   4
C3H5OO                  C   3H   5O   2     G    300.00   3500.00 1800.00      1
 7.69230110e+00 2.05361077e-02-9.61589847e-06 2.15332094e-09-1.88909485e-13    2
 6.21484234e+03-1.04053755e+01 2.96424215e+00 3.10429054e-02-1.83715632e-05    3
 5.39615972e-09-6.39303761e-13 7.91694356e+03 1.51838658e+01                   4
C3H5OOH                 C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.21377197e+01 1.68585481e-02-6.94275126e-06 1.36958900e-09-1.07427460e-13    2
-1.25265904e+04-3.57194708e+01 2.24651097e+00 3.88390118e-02-2.52598044e-05    3
 8.15368275e-09-1.04966270e-12-8.96575529e+03 1.78138141e+01                   4
C3H6                    C   3H   6          G    300.00   3500.00 1800.00      1
 9.21549195e+00 1.10096151e-02-2.72165887e-06 1.69301120e-10 1.25058839e-14    2
-2.15028535e+03-2.75773224e+01-2.61886761e-01 3.20704567e-02-2.02723602e-05    3
 6.66956086e-09-8.90307969e-13 1.26157099e+03 2.37162283e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1720.00      1
 6.42754902e+00 2.00818525e-02-6.55464685e-06 4.84306793e-10 5.68893699e-14    2
-1.48035725e+04-9.71995026e+00-9.99780843e-02 3.52621481e-02-1.97932767e-05    3
 5.61555868e-09-6.88932126e-13-1.25581031e+04 2.53116313e+01                   4
C3H6O2                  C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.08721654e+01 1.63593216e-02-6.08637842e-06 1.10130850e-09-8.02911326e-14    2
-4.55272952e+04-2.70748520e+01 2.66105929e+00 3.46062241e-02-2.12921305e-05    3
 6.73306853e-09-8.62480026e-13-4.25712970e+04 1.73653673e+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   3500.00  700.00      1
-9.77279434e-01 5.24983747e-02-3.09762338e-05 8.32680251e-09-8.38156520e-13    2
-2.70767712e+04 3.27194912e+01 3.71554492e+00 2.56822356e-02 2.64869216e-05    3
-4.64000121e-08 1.87071344e-11-2.77337666e+04 1.17531393e+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   3500.00 1670.00      1
 1.20273024e+01 2.23669330e-02-9.25510611e-06 1.83134653e-09-1.43510571e-13    2
-2.87878078e+04-3.43698022e+01 1.14029559e+00 4.84435961e-02-3.26772586e-05    3
 1.11815072e-08-1.54323522e-12-2.51515476e+04 2.37368269e+01                   4
C3H8                    C   3H   8          G    300.00   3500.00 1800.00      1
 1.08596364e+01 1.35766563e-02-3.19926248e-06 1.41615801e-10 2.35898562e-14    2
-1.80884704e+04-3.69486914e+01-1.25512725e+00 4.04983533e-02-2.56340099e-05    3
 8.45078153e-09-1.13046094e-12-1.37271555e+04 2.86189366e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00 1050.00      1
 8.50275797e+00 6.97445022e-03-2.53297106e-06 4.33287765e-10-2.93611469e-14    2
 5.31727553e+04-2.08807943e+01 2.90907865e+00 2.82837048e-02-3.29747633e-05    3
 1.97614098e-08-4.63129497e-12 5.43474279e+04 6.37839155e+00                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590365e-03 1.80568199e-06-9.30237202e-10 1.18077197e-13    2
 6.01811751e+04-4.25791500e+01 2.34662667e+00 2.83894138e-02-2.35278181e-05    3
 9.69177542e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H3O                   C   4H   3O   1     G    300.00   3500.00 1240.00      1
 8.44125905e+00 1.62911136e-02-8.34126436e-06 2.01436766e-09-1.87394603e-13    2
 1.94535776e+04-2.27855078e+01-5.90872253e+00 6.25813767e-02-6.43375505e-05    3
 3.21198978e-08-6.25705794e-12 2.30123730e+04 4.95317026e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1190.00      1
 6.36293592e+00 1.66610000e-02-7.54220850e-06 1.59521425e-09-1.28415834e-13    2
 3.13137240e+04-8.19255288e+00 4.03184847e-01 3.66937767e-02-3.27936077e-05    3
 1.57416564e-08-3.10035746e-12 3.27321448e+04 2.15965194e+01                   4
C4H4O                   C   4H   4O   1     G    300.00   3500.00 1250.00      1
 8.37486466e+00 1.95634451e-02-9.90167121e-06 2.37694382e-09-2.20517698e-13    2
-9.41817580e+03-2.52053384e+01-7.59507781e+00 7.06672610e-02-7.12262503e-05    3
 3.50833860e-08-6.76180613e-12-5.42569018e+03 5.54039922e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794385e-03 4.88814513e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742307e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H6                    C   4H   6          G    300.00   3500.00 1550.00      1
 9.55395345e+00 1.51364811e-02-4.78509457e-06 6.14955374e-10-2.23809938e-14    2
 8.63284693e+03-2.77966685e+01-1.04533857e+00 4.24894928e-02-3.12557510e-05    3
 1.20001840e-08-1.85870818e-12 1.19186275e+04 2.79839806e+01                   4
C4H6O2                  C   4H   6O   2     G    300.00   3500.00 1800.00      1
 7.01919581e+00 2.89919962e-02-1.39811163e-05 3.22750474e-09-2.90888810e-13    2
-4.36055710e+04-7.47846940e+00 9.15158242e-01 4.25565241e-02-2.52848896e-05    3
 7.41408744e-09-8.72358628e-13-4.14081175e+04 2.55578553e+01                   4
C4H7OH                  C   4H   8O   1     G    300.00   3500.00 1460.00      1
 1.00981665e+01 2.15734935e-02-6.74008418e-06 9.16825971e-10-4.16200161e-14    2
-2.37290909e+04-2.45741592e+01-2.55531336e-01 4.99397889e-02-3.58835384e-05    3
 1.42243393e-08-2.32030381e-12-2.07058111e+04 2.92946643e+01                   4
C4H8O                   C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.12815996e+01 2.48463701e-02-1.13234700e-05 2.47069946e-09-2.12413507e-13    2
-2.03756688e+04-3.84267373e+01-2.94845122e+00 5.64687053e-02-3.76754160e-05    3
 1.22306795e-08-1.56796629e-12-1.52528505e+04 3.85892666e+01                   4
C4H9CHO                 C   5H  10O   1     G    300.00   3500.00  760.00      1
-1.78433179e+00 6.31204386e-02-3.60836198e-05 9.48321920e-09-9.39522544e-13    2
-2.97113508e+04 3.92478712e+01 5.53299014e+00 2.46082180e-02 3.99273421e-05    3
-5.71930632e-08 2.09934651e-11-3.08235837e+04 5.95416540e+00                   4
C4H9OOH                 C   4H  10O   2     G    300.00   3500.00 1780.00      1
 1.73966948e+01 2.30088698e-02-8.34646932e-06 1.39883190e-09-9.01677555e-14    2
-3.38614042e+04-6.23628946e+01 1.12895120e+00 5.95655969e-02-3.91527000e-05    3
 1.29367460e-08-1.71066131e-12-2.80700874e+04 2.54997628e+01                   4
C5EN-OO                 C   5H   9O   2     G    300.00   3500.00 1280.00      1
 1.00840321e+01 3.69913036e-02-1.74216180e-05 3.93130749e-09-3.47257402e-13    2
-8.98415155e+02-1.96513637e+01 4.09897281e-01 6.72229749e-02-5.28493577e-05    3
 2.23832553e-08-3.95115346e-12 1.57816336e+03 2.94089022e+01                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   3500.00 1160.00      1
 1.36699765e+01 4.21231935e-02-2.15503712e-05 5.21806336e-09-4.87293014e-13    2
-1.42354804e+04-3.35883364e+01 5.24578583e-01 8.74521518e-02-8.01654035e-05    3
 3.89048635e-08-7.74737926e-12-1.11857480e+04 3.17816498e+01                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   3500.00 1580.00      1
 1.69833146e+01 2.73095032e-02-1.19226853e-05 2.48166925e-09-2.03420392e-13    2
-3.51234520e+04-5.58041780e+01 1.44561329e+00 6.66454559e-02-4.92669442e-05    3
 1.82387405e-08-2.69662788e-12-3.02135384e+04 2.62635800e+01                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   3500.00 1420.00      1
 1.28791275e+01 3.32930454e-02-1.55378924e-05 3.46674396e-09-3.02869803e-13    2
 3.23011716e+03-3.38507184e+01 1.34404411e+00 6.57862381e-02-4.98616876e-05    3
 1.95812018e-08-3.13992224e-12 6.50608085e+03 2.58442475e+01                   4
C5H4O2                  C   5H   4O   2     G    300.00   3500.00 1430.00      1
 1.05158962e+01 2.23224229e-02-1.09267096e-05 2.56683236e-09-2.34844997e-13    2
-2.33303219e+04-2.94000374e+01-1.81996644e+00 5.68283325e-02-4.71217197e-05    3
 1.94409629e-08-3.18486782e-12-1.98022652e+04 3.45255921e+01                   4
C5H5O                   C   5H   5O   1     G    300.00   3500.00 1450.00      1
 1.05801390e+01 2.13128784e-02-9.63052935e-06 2.09384798e-09-1.79321204e-13    2
 1.62543411e+04-3.26154734e+01-4.01979397e+00 6.15885556e-02-5.12950230e-05    3
 2.12499370e-08-3.48209517e-12 2.04883217e+04 4.32455666e+01                   4
C5H7                    C   5H   7          G    300.00   3500.00 1430.00      1
 7.72404525e+00 2.56072196e-02-8.76350316e-06 8.66193959e-10 3.30416650e-14    2
 2.30808142e+04-1.69352935e+01 2.31765047e-01 4.65646468e-02-3.07468184e-05    3
 1.11148258e-08-1.75867718e-12 2.52236063e+04 2.18904247e+01                   4
C5H8                    C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829159e+00 2.51033002e-02-8.43679234e-06 8.19905621e-10 3.11426511e-14    2
 4.67953300e+03-2.40439628e+01 1.19183502e+00 4.68276543e-02-3.12245763e-05    3
 1.14435811e-08-1.82614328e-12 6.90073958e+03 1.62025638e+01                   4
C5H8O                   C   5H   8O   1     G    300.00   3500.00 1330.00      1
 6.70800688e+00 3.65243775e-02-1.77765821e-05 4.15639148e-09-3.79163309e-13    2
-5.52771782e+03-9.67918417e+00-5.12640161e+00 7.21165834e-02-5.79181678e-05    3
 2.42774871e-08-4.16132413e-12-2.37976516e+03 5.07899199e+01                   4
C5H8O4                  C   5H   8O   4     G    300.00   3500.00 1230.00      1
 1.19601536e+01 3.99450843e-02-1.95947373e-05 4.60940117e-09-4.22302290e-13    2
-8.26385858e+04-2.91875208e+01-6.95683231e+00 1.01463738e-01-9.46174851e-05    3
 4.52721371e-08-8.68708602e-12-7.79850073e+04 6.59920851e+01                   4
C5H9CHO                 C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.08416239e+01 4.20296686e-02-2.00742994e-05 4.57927363e-09-4.08519043e-13    2
-3.59631714e+04-3.80017802e+01-6.51363638e+00 8.05969136e-02-5.22136702e-05    3
 1.64827443e-08-2.06177886e-12-2.97152777e+04 5.59285088e+01                   4
C6H10O5                 C   6H  10O   5     G    300.00   3500.00 1220.00      1
 1.54889718e+01 4.96354387e-02-2.45944509e-05 5.82332585e-09-5.35665863e-13    2
-1.09180509e+05-4.81819837e+01-7.95116461e+00 1.26488345e-01-1.19085729e-04    3
 5.74579042e-08-1.11165221e-11-1.03461116e+05 6.95642163e+01                   4
C6H2                    C   6H   2          G    300.00   3500.00 1100.00      1
 1.20007067e+01 9.35747205e-03-3.45039279e-06 5.96931921e-10-4.08067421e-14    2
 8.10797696e+04-3.61630610e+01 4.40206371e+00 3.69889013e-02-4.11296144e-05    3
 2.34328238e-08-5.23078218e-12 8.27514710e+04 1.22022725e+00                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194523e+01 1.16137832e-02-4.19264523e-06 6.84693072e-10-4.17887568e-14    2
 8.26280760e+04-3.29876543e+01 4.46601450e+00 3.41999583e-02-2.98587533e-05    3
 1.36473739e-08-2.49684195e-12 8.45957836e+04 5.04018537e+00                   4
C6H4                    C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447675e+01 6.21306708e-03-9.80963858e-07 8.00594635e-11-2.88320770e-15    2
 5.49568894e+04-6.59208082e+01-1.17305610e+00 6.09713718e-02-6.13761529e-05    3
 2.96855443e-08-5.44506791e-12 6.00209374e+04 2.96241244e+01                   4
C6H4C2H                 C   8H   5          G    300.00   3500.00 1490.00      1
 3.21415686e+01-1.98168404e-02 2.64282529e-05-1.09843473e-08 1.50630597e-12    2
 5.44964091e+04-1.47026437e+02-4.78252619e+00 7.93082463e-02-7.33621030e-05    3
 3.36645815e-08-5.98512503e-12 6.54997893e+04 4.58354239e+01                   4
C6H4CH3                 C   7H   7          G    300.00   3500.00 1450.00      1
 1.23344954e+01 2.38147082e-02-7.01721971e-06 3.58622104e-10 7.92842393e-14    2
 2.97091697e+04-3.94240761e+01-4.14387803e+00 6.92722902e-02-5.40423045e-05    3
 2.19793508e-08-3.64842760e-12 3.44878980e+04 4.61973136e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929577e+01 1.29021286e-02-2.02976642e-06-3.72417846e-10 8.59745727e-14    2
-2.22100459e+04-6.49015838e+01-5.23446578e+00 7.73770890e-02-7.06201498e-05    3
 3.20580235e-08-5.66410367e-12-1.58009124e+04 5.25540058e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1690.00      1
 2.37494889e+01-3.74826288e-03 7.22829016e-06-2.69927706e-09 3.10032681e-13    2
 2.93571719e+04-1.07010346e+02-4.30972117e+00 6.26640688e-02-5.17175663e-05    3
 2.05535263e-08-3.12973113e-12 3.88411849e+04 4.30825907e+01                   4
C6H5C2H                 C   8H   6          G    300.00   3500.00 1330.00      1
 1.36301627e+01 2.67826138e-02-1.18276978e-05 2.56807250e-09-2.21616638e-13    2
 3.04381476e+04-4.83434869e+01-3.73085925e+00 7.89962135e-02-7.07152163e-05    3
 3.20856256e-08-5.77002888e-12 3.50561794e+04 4.03644060e+01                   4
C6H5C2H2                C   8H   7          G    300.00   3500.00 1690.00      1
 1.77155600e+01 2.19043174e-02-8.07391246e-06 1.39474201e-09-9.41524347e-14    2
 3.81394494e+04-7.01114193e+01-2.50848763e+00 6.97718858e-02-5.05599199e-05    3
 1.81545083e-08-2.57340780e-12 4.49751775e+04 3.80700548e+01                   4
C6H5C2H3                C   8H   8          G    300.00   3500.00 1420.00      1
 1.57612121e+01 2.51344730e-02-7.08348959e-06 3.12355848e-10 8.22985790e-14    2
 1.01346894e+04-5.95859946e+01-4.61890423e+00 8.25432514e-02-6.77265654e-05    3
 2.87832834e-08-4.93018867e-12 1.59226425e+04 4.58827137e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1440.00      1
 2.29999925e+01 5.23551496e-02-1.62023052e-05 1.06346924e-09 1.48747565e-13    2
 3.20131872e+03-9.18704227e+01-1.05589612e+01 1.45574466e-01-1.13305759e-04    3
 4.60187721e-08-7.65599251e-12 1.28662974e+04 8.22691715e+01                   4
C6H5C2H5                C   8H  10          G    300.00   3500.00 1440.00      1
 1.53992430e+01 3.11284429e-02-9.32920034e-06 5.29654938e-10 9.71609974e-14    2
-4.32725762e+03-5.77491740e+01-6.11786341e+00 9.08981829e-02-7.15893461e-05    3
 2.93537965e-08-4.90703025e-12 1.86966902e+03 5.39044909e+01                   4
C6H5CH2C6H5             C  13H  12          G    300.00   3500.00 1440.00      1
 2.36600260e+01 4.20961068e-02-1.18756749e-05 4.02369975e-10 1.68531444e-13    2
 4.50897730e+03-9.76688099e+01-1.18613481e+01 1.40766591e-01-1.14657429e-04    3
 4.79865153e-08-8.09260490e-12 1.47391331e+04 8.66539117e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799879e-06 4.38368241e-10 8.64078959e-14    2
-1.87828963e+04-3.81332333e+01-6.02884975e+00 7.77532977e-02-6.10481840e-05    3
 2.48568442e-08-4.12367417e-12-1.33857950e+04 5.85676633e+01                   4
C6H5CHO                 C   7H   6O   1     G    300.00   3500.00 1770.00      1
 2.73588480e+01 2.45725463e-03 5.41130341e-06-2.58531717e-09 3.21649872e-13    2
-1.76429542e+04-1.23608292e+02-6.55705980e+00 7.91033740e-02-5.95430351e-05    3
 2.18795937e-08-3.13384602e-12-5.63672287e+03 5.93816475e+01                   4
C6H5O                   C   6H   5O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658729e-02-6.67332779e-06 1.12237517e-09-7.10809502e-14    2
 4.07683820e+02-4.72500520e+01-4.80707078e+00 7.32685627e-02-6.95172935e-05    3
 3.28617518e-08-6.08232652e-12 5.22565416e+03 4.58618544e+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   3500.00 1380.00      1
 1.25085136e+01 3.49906122e-02-1.63096082e-05 3.64836832e-09-3.19988393e-13    2
-1.52038795e+04-4.20406499e+01-5.29461551e+00 8.65938851e-02-7.24001222e-05    3
 3.07452350e-08-5.22884105e-12-1.02902159e+04 4.95832512e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867712e+01 2.02277643e-02-7.36599500e-06 1.21196288e-09-7.46105018e-14    2
-1.80542263e+04-5.08485811e+01-5.47325435e+00 7.87541571e-02-7.33732049e-05    3
 3.42982836e-08-6.29384372e-12-1.28778595e+04 4.85843830e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1550.00      1
 1.57365829e+01 1.24444139e-02-2.08242468e-06-1.90555168e-10 5.60938650e-14    2
 2.37538837e+03-6.60380946e+01-6.33361145e+00 6.93997541e-02-5.72004958e-05    3
 2.35161421e-08-3.76756698e-12 9.21714860e+03 5.01102066e+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   3500.00 1770.00      1
 1.98638073e+01 1.79335016e-02-5.95408859e-06 8.93593939e-10-4.95459880e-14    2
-4.95264845e+04-7.44496694e+01 7.10718582e-01 6.12173180e-02-4.26352889e-05    3
 1.47094886e-08-2.00094354e-12-4.27462910e+04 2.88889342e+01                   4
C6H8O4                  C   6H   8O   4     G    300.00   3500.00 1300.00      1
 1.58073709e+01 3.77998882e-02-1.77241312e-05 3.97560136e-09-3.49009860e-13    2
-7.78788467e+04-5.15128322e+01-4.55493836e+00 1.00453147e-01-9.00163533e-05    3
 4.10485358e-08-7.47842033e-12-7.25846463e+04 5.20658817e+01                   4
C7DIONE                 C   7H  12O   2     G    300.00   3500.00  700.00      1
-7.55853587e-01 8.24536116e-02-4.58824665e-05 1.18274999e-08-1.15807940e-12    2
-3.67546790e+04 2.64722477e+01 3.52180397e+00 5.80098541e-02 6.49701379e-06    3
-3.80577194e-08 1.66580704e-11-3.73535510e+04 7.36075600e+00                   4
C7H15COCHO              C   9H  16O   2     G    300.00   3500.00 1780.00      1
 3.02050983e+01 3.84107591e-02-1.30454122e-05 2.02881682e-09-1.19348346e-13    2
-6.67956450e+04-1.25747051e+02 3.59041588e-01 1.05480549e-01-6.95648985e-05    3
 2.31971638e-08-3.09243078e-12-5.61704488e+04 3.54525548e+01                   4
C7H7                    C   7H   7          G    300.00   3500.00 1450.00      1
 1.55564029e+01 1.97467971e-02-4.90102499e-06-1.06746050e-11 9.16513058e-14    2
 1.67098727e+04-6.15086686e+01-4.40172355e+00 7.48036976e-02-6.18564392e-05    3
 2.61757227e-08-4.42324479e-12 2.24977294e+04 4.21934668e+01                   4
C7H8                    C   7H   8          G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799879e-06 4.38368241e-10 8.64078959e-14    2
-5.64471283e+02-4.45247833e+01-6.02884975e+00 7.77532977e-02-6.10481840e-05    3
 2.48568442e-08-4.12367417e-12 4.83263000e+03 5.21761133e+01                   4
C7KETONE                C   7H  14O   1     G    300.00   3500.00 1800.00      1
 1.82994273e+01 4.14393597e-02-1.71834162e-05 3.42714287e-09-2.72037363e-13    2
-4.27848802e+04-6.59785823e+01-2.29236271e-01 8.26141675e-02-5.14957561e-05    3
 1.61354169e-08-2.03707542e-12-3.61145614e+04 3.43024100e+01                   4
C8H10O3                 C   8H  10O   3     G    300.00   3500.00 1280.00      1
 2.98957517e+01 4.73870505e-02-2.11603212e-05 4.60350399e-09-3.96349099e-13    2
-7.02119467e+04-1.21160681e+02-3.09348688e+00 1.50478421e-01-1.41970521e-04    3
 6.75254832e-08-1.26857982e-11-6.17667016e+04 4.61370519e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874492e-03-2.93037080e-06 2.89537341e-10 2.52405898e-16    2
 1.07885460e+05-5.89733614e+01 1.87361722e-01 7.06952484e-02-8.88216494e-05    3
 5.43092094e-08-1.27402363e-11 1.11295389e+05 1.95626382e+01                   4
C8H9                    C   8H   9          G    300.00   3500.00 1570.00      1
 2.45973914e+01 1.20503967e-02 5.66754133e-07-1.10955314e-09 1.57308310e-13    2
 1.65948730e+04-1.06442126e+02-5.12604623e+00 8.77789001e-02-7.17853192e-05    3
 2.96131956e-08-4.73484913e-12 2.59280324e+04 5.03637968e+01                   4
C9H10O2                 C   9H  10O   2     G    300.00   3500.00 1620.00      1
 2.64048781e+01 2.84903123e-02-1.03289369e-05 1.78607618e-09-1.22280426e-13    2
-3.71439509e+04-1.10770565e+02-2.04331024e+00 9.87327525e-02-7.53682334e-05    3
 2.85512188e-08-4.25270367e-12-2.79267379e+04 4.01996488e+01                   4
CH                      C   1H   1          G    300.00   3500.00 1720.00      1
 1.56762354e+00 3.35441204e-03-1.29971595e-06 2.40500907e-10-1.78141164e-14    2
 7.11686733e+04 1.27712404e+01 3.85901271e+00-1.97439999e-03 3.34750385e-06    3
-1.56074708e-09 2.43995183e-13 7.03804355e+04 4.73936215e-01                   4
CH2                     C   1H   2          G    300.00   3500.00  900.00      1
 3.24505871e+00 2.75395076e-03-7.68471343e-07 8.23040037e-11-1.89900250e-15    2
 4.54794580e+04 4.28187007e+00 3.99717917e+00-5.88806826e-04 4.80279129e-06    3
-4.04455721e-09 1.14445133e-12 4.53440763e+04 7.32567433e-01                   4
CH2C3H5                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075606e-06 3.82147973e-10 5.73994806e-14    2
 1.98988324e+04-1.80212793e+01-3.29329051e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
CH2CCH3                 C   3H   5          G    300.00   3500.00 1800.00      1
 1.00124373e+01 7.55815802e-03-1.17096962e-06-2.01794819e-10 4.72987983e-14    2
 2.78641947e+04-2.75169832e+01 6.10512020e-01 2.84513252e-02-1.85819423e-05    3
 6.24671358e-09-8.48327368e-13 3.12488878e+04 2.33681976e+01                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   3500.00 1590.00      1
 1.05858550e+01 1.29956017e-02-4.76361255e-06 7.49449815e-10-3.96847802e-14    2
 3.10513348e+03-2.93262371e+01 1.05972039e+00 3.69607201e-02-2.73722149e-05    3
 1.02289476e-08-1.53017186e-12 6.13444428e+03 2.10494483e+01                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.17572858e+01 2.41574264e-02-9.72976868e-06 1.89143875e-09-1.46945289e-13    2
-1.45672160e+04-3.14377946e+01 8.93764133e-01 4.82985857e-02-2.98474014e-05    3
 9.34241382e-09-1.18180294e-12-1.06563482e+04 2.73578508e+01                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.49770379e+00 1.77061096e-02-6.68456978e-06 1.20981994e-09-8.73179586e-14    2
-1.07976200e+04-2.07829255e+01 1.04629052e+00 3.64870279e-02-2.23353351e-05    3
 7.00639969e-09-8.92398479e-13-7.75511123e+03 2.49578861e+01                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097165e-06 1.27900113e-09-8.37238502e-14    2
-1.74897435e+04-4.46134901e+01 9.11733056e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH2CHCH2                C   3H   5          G    300.00   3500.00 1800.00      1
 1.31270112e+01 3.37812631e-03 1.30787951e-06-8.72502093e-10 1.13779857e-13    2
 1.38569110e+04-4.71985703e+01 1.45788193e-01 3.22252886e-02-2.27314224e-05    3
 8.03094306e-09-1.12280975e-12 1.85301513e+04 2.30585168e+01                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   3500.00 1780.00      1
 1.38129918e+01 2.02819032e-02-7.03372780e-06 1.12439860e-09-6.86002896e-14    2
-1.64045579e+04-4.42517079e+01 2.32452600e-01 5.07999690e-02-3.27511989e-05    3
 1.07564103e-08-1.42141092e-12-1.15698860e+04 2.90972641e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1030.00      1
 3.66502520e+00 1.44768244e-02-7.23266377e-06 1.70580456e-09-1.56345856e-13    2
-3.68579193e+01 5.92341850e+00 2.15742069e-01 2.78720987e-02-2.67403448e-05    3
 1.43321353e-08-3.22098924e-12 6.73694406e+02 2.26661724e+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   3500.00 1380.00      1
 6.32694430e+00 2.38762490e-02-1.07376178e-05 2.33737032e-09-2.01069469e-13    2
-1.14217376e+04-3.95690500e+00 6.40756935e-01 4.03579515e-02-2.86525118e-05    3
 1.09919085e-08-1.76892059e-12-9.85234986e+03 2.53070892e+01                   4
CH2CHOOHCHO             C   3H   5O   3     G    300.00   3500.00 1300.00      1
 1.09154411e+01 2.11069264e-02-1.04347901e-05 2.43633157e-09-2.20224944e-13    2
-1.35446352e+04-2.42468452e+01 1.81101363e+00 4.91205495e-02-4.27582013e-05    3
 1.90124399e-08-3.40793808e-12-1.11774841e+04 2.20654311e+01                   4
CH2CN                   C   2H   2N   1     G    300.00   3500.00  980.00      1
 4.41880974e+00 9.83430327e-03-4.98991807e-06 1.22319871e-09-1.17396557e-13    2
 2.92390343e+04 2.02769260e+00 2.71162977e+00 1.68023848e-02-1.56553489e-05    3
 8.47859386e-09-1.96826267e-12 2.95736416e+04 1.02293594e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1410.00      1
 6.03578795e+00 5.81722422e-03-1.93206512e-06 2.83140054e-10-1.50051612e-14    2
-8.58422380e+03-7.64505060e+00 2.49197065e+00 1.58706066e-02-1.26271528e-05    3
 5.33991909e-09-9.11597189e-13-7.58486732e+03 1.06694385e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  930.00      1
 1.06639253e+00 1.06960337e-02-5.54447373e-06 1.36053696e-09-1.28442554e-13    2
-1.46324373e+04 1.74071779e+01 3.13463322e+00 1.80037482e-03 8.80336316e-06    3
-8.92465077e-09 2.63639286e-12-1.50171301e+04 7.57920580e+00                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1590.00      1
 7.61004151e+00 1.40239019e-03 1.05265418e-06-5.61972284e-10 7.11209072e-14    2
-5.04985629e+03-1.55757586e+01 1.95857131e+00 1.56199253e-02-1.23601148e-05    3
 5.06183022e-09-8.13124769e-13-3.25268877e+03 1.43100973e+01                   4
CH2OOCH2CHO             C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.06998539e+01 2.42793089e-02-1.34097218e-05 3.42673974e-09-3.32159552e-13    2
-2.14126656e+04-2.48508794e+01 2.93009251e+00 4.15454454e-02-2.77981689e-05    3
 8.75579421e-09-1.07230601e-12-1.86155515e+04 1.72006902e+01                   4
CH2OOCHOOHCHO           C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549192e+01 1.08256409e-02-3.75393277e-06 5.88014009e-10-3.47282962e-14    2
-3.59900210e+04-7.93559883e+01 5.41191662e+00 4.64767576e-02-3.34631967e-05    3
 1.15914451e-08-1.56298261e-12-3.02145401e+04 7.47208818e+00                   4
CH2OOHCHCHO             C   3H   5O   3     G    300.00   3500.00  700.00      1
 1.84816700e+00 3.99042619e-02-2.38947704e-05 6.48850081e-09-6.57628290e-13    2
-1.48991977e+04 2.15340498e+01 5.44326670e+00 1.93608350e-02 2.01268587e-05    3
-3.54368602e-08 1.43157149e-11-1.54025117e+04 5.47205385e+00                   4
CH2OOHCHOOCHO           C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549192e+01 1.08256409e-02-3.75393277e-06 5.88014009e-10-3.47282962e-14    2
-3.59900210e+04-7.93559883e+01 5.41191662e+00 4.64767576e-02-3.34631967e-05    3
 1.15914451e-08-1.56298261e-12-3.02145401e+04 7.47208818e+00                   4
CH2S                    C   1H   2          G    300.00   3500.00  900.00      1
 2.57518275e+00 4.11179659e-03-1.68232435e-06 3.44404948e-10-2.93085968e-14    2
 5.01958500e+04 6.99914504e+00 4.62572654e+00-5.00173140e-03 1.35068890e-05    3
-1.09068642e-08 3.09604394e-12 4.98267521e+04-2.67749711e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1270.00      1
 2.57723974e+00 6.62601164e-03-2.54906392e-06 4.67320141e-10-3.34867663e-14    2
 1.65488693e+04 6.94195966e+00 3.53327401e+00 3.61488008e-03 1.00739068e-06    3
-1.39958516e-09 3.34014277e-13 1.63060366e+04 2.10113860e+00                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936624e+01 3.24954978e-02-1.30480618e-05 2.52260906e-09-1.95492396e-13    2
-2.87396993e+03-1.14905139e+02-1.85059487e+00 9.45938472e-02-6.47966864e-05    3
 2.16887663e-08-2.85745868e-12 7.18596268e+03 3.63350107e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191869e+01 2.86451308e-02-9.80098219e-06 1.51374083e-09-8.72237944e-14    2
-2.13626711e+04-1.32660114e+02-1.76841814e+00 9.72842531e-02-6.70002508e-05    3
 2.26986551e-08-3.02957300e-12-1.02431333e+04 3.45100483e+01                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   3500.00  700.00      1
 2.02076663e+00 4.09903683e-02-2.06486866e-05 5.00507647e-09-4.71523451e-13    2
-1.40718373e+04 2.15880986e+01 3.53447938e+00 3.23405812e-02-2.11342851e-06    3
-1.26475503e-08 5.83298611e-12-1.42837571e+04 1.48252130e+01                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.16093380e+01 2.56981798e-02-1.09676558e-05 2.25993093e-09-1.85313976e-13    2
-1.31948148e+04-3.43573902e+01 5.90549372e-02 5.13654755e-02-3.23570689e-05    3
 1.01819358e-08-1.28559243e-12-9.03671291e+03 2.81551514e+01                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.30151659e+01 2.21750012e-02-8.49156594e-06 1.54860371e-09-1.12013678e-13    2
-1.79081220e+04-4.01994427e+01 1.75489331e+00 4.71978292e-02-2.93439226e-05    3
 9.27169878e-09-1.18466577e-12-1.38544238e+04 2.07435017e+01                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.07749584e+00 1.96975457e-02-8.18089073e-06 1.64328968e-09-1.31786153e-13    2
-9.31061125e+03-2.21687275e+01 2.91958855e-01 3.92209612e-02-2.44504037e-05    3
 7.66903521e-09-9.68695255e-13-6.14781793e+03 2.53804314e+01                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.15124775e+01 2.41072597e-02-9.86401997e-06 1.98674692e-09-1.62119892e-13    2
-1.58991633e+04-3.03580006e+01 1.53457350e-01 4.93495266e-02-3.08992425e-05    3
 9.77757006e-09-1.24417866e-12-1.18099160e+04 3.11193861e+01                   4
CH3CH2CHOCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.30434362e+01 2.38164771e-02-9.82552432e-06 1.93897534e-09-1.51918988e-13    2
-1.58538336e+04-4.35088383e+01 4.17731726e-02 5.27090615e-02-3.39026780e-05    3
 1.08564397e-08-1.39045570e-12-1.11732349e+04 2.68588742e+01                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   3500.00 1620.00      1
 8.28181025e+00 2.00744959e-02-8.21041648e-06 1.62349331e-09-1.27917758e-13    2
-1.30492834e+04-1.56179098e+01 1.73835403e+00 3.62311779e-02-2.31703072e-05    3
 7.77982697e-09-1.07796925e-12-1.09292035e+04 1.91072184e+01                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097165e-06 1.27900113e-09-8.37238502e-14    2
-1.74897435e+04-4.46134901e+01 9.11733056e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   3500.00 1430.00      1
 8.72382272e+00 3.04342830e-02-1.39185549e-05 3.06043861e-09-2.64689231e-13    2
-1.80661273e+04-1.71435098e+01 1.27395834e+00 5.12730645e-02-3.57774166e-05    3
 1.32510501e-08-2.04626467e-12-1.59354661e+04 2.14624055e+01                   4
CH3CH3-C5H6             C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755546e+01 3.27318283e-02-1.05955708e-05 1.52102630e-09-7.69415914e-14    2
-6.19682930e+03-5.37226046e+01-1.29247813e+00 8.36265847e-02-6.88720094e-05    3
 3.11782470e-08-5.73671653e-12-1.82980473e+03 3.11918393e+01                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.15124775e+01 2.41072597e-02-9.86401997e-06 1.98674692e-09-1.62119892e-13    2
-1.58991633e+04-3.03580006e+01 1.53457350e-01 4.93495266e-02-3.08992425e-05    3
 9.77757006e-09-1.24417866e-12-1.18099160e+04 3.11193861e+01                   4
CH3CHCH2OCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.38488385e+01 2.14834842e-02-8.03028843e-06 1.42167056e-09-9.95437051e-14    2
-1.51249440e+04-4.82209549e+01-4.69026374e-01 5.33009618e-02-3.45448531e-05    3
 1.12418797e-08-1.46346164e-12-9.97051265e+03 2.92703168e+01                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 7.64501934e+00 2.06996931e-02-8.77824684e-06 1.84245353e-09-1.55992331e-13    2
-1.15050426e+04-1.08131884e+01 5.39035202e-01 3.64907690e-02-2.19374767e-05    3
 6.71624238e-09-8.32907449e-13-8.94688828e+03 2.76458802e+01                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   3500.00 1450.00      1
 8.91411879e+00 2.94184843e-02-1.30488503e-05 2.81020956e-09-2.39749810e-13    2
-1.71145335e+04-1.85255698e+01 6.16106328e-01 5.23095531e-02-3.67292664e-05    3
 1.36977572e-08-2.11691319e-12-1.47081099e+04 2.45907827e+01                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.11524016e+01 2.52912378e-02-1.05179486e-05 2.12392650e-09-1.71553011e-13    2
-1.78095410e+04-2.94209720e+01 6.76902371e-01 4.85701251e-02-2.99170213e-05    3
 9.30876825e-09-1.16944770e-12-1.40383613e+04 2.72746153e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.27018126e+00 1.06201871e-02-3.82264672e-06 6.56340789e-10-4.60549581e-14    2
-2.29794782e+04-8.60119259e+00 9.91751377e-01 2.23500313e-02-1.35975169e-05    3
 4.27666307e-09-5.48877497e-13-2.10792434e+04 1.99667711e+01                   4
CH3CHOH                 C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.00303702e+00 2.30237358e-02-1.19372743e-05 2.98274467e-09-2.88183748e-13    2
-6.17751011e+03 2.39401608e+01 1.83915526e+00 1.82459173e-02-1.69909177e-06    3
-6.76790535e-09 3.19419126e-12-6.29456667e+03 2.02045961e+01                   4
CH3CHOOCHO              C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.58771657e+01 1.28699615e-02-5.29703385e-06 1.04001953e-09-8.12487153e-14    2
-2.38887629e+04-5.44666587e+01 3.38301196e+00 4.06347476e-02-2.84343556e-05    3
 9.60939795e-09-1.27144016e-12-1.93908676e+04 1.31543077e+01                   4
CH3CN                   C   2H   3N   1     G    300.00   3500.00  700.00      1
 2.02660925e+00 1.64402545e-02-8.54290907e-06 2.13740318e-09-2.08581596e-13    2
 8.61823027e+03 1.31030643e+01 2.36621609e+00 1.44996440e-02-4.38445795e-06    3
-1.82302645e-09 1.20585756e-12 8.57068531e+03 1.15857868e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 5.59449005e+00 8.95063669e-03-3.42706569e-06 6.39554414e-10-4.91680987e-14    2
-5.31931220e+03-3.46466160e+00 1.83189171e+00 1.73119663e-02-1.03948404e-05    3
 3.22021171e-09-4.07592723e-13-3.96477680e+03 1.68993055e+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483421e-03 1.65900438e-06-8.55133987e-10 9.82287242e-14    2
-2.73756816e+04-4.36816972e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1760.00      1
 1.54960865e+01 1.58758106e-03 2.24425901e-06-9.74237206e-10 1.03773065e-13    2
-4.69655432e+04-5.18401164e+01 3.62388957e+00 2.85698467e-02-2.07519902e-05    3
 7.73646324e-09-1.13354234e-12-4.27865299e+04 1.21478877e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 9.24187097e+00 1.34946785e-02-5.23722666e-06 9.72748882e-10-7.19834442e-14    2
-8.04571079e+03-2.24258259e+01 1.82620860e+00 2.99739283e-02-1.89699348e-05    3
 6.05893707e-09-7.78398470e-13-5.37607233e+03 1.77092859e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00  700.00      1
 8.22157368e-01 3.18964631e-02-1.68324056e-05 4.20706053e-09-4.04124926e-13    2
-2.74737271e+04 2.17873546e+01 1.03654018e+00 3.06714184e-02-1.42073099e-05    3
 1.70696939e-09 4.88764769e-13-2.75037407e+04 2.08295464e+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   3500.00 1270.00      1
 6.71652579e+00 2.35306498e-02-1.06144747e-05 2.31761627e-09-1.99886320e-13    2
-1.44175086e+04-7.90476332e+00 1.21649821e+00 4.08535713e-02-3.10746182e-05    3
 1.30578491e-08-2.31410538e-12-1.30205016e+04 1.99442900e+01                   4
CH3COOH                 C   2H   4O   2     G    300.00   3500.00 1410.00      1
 7.83491620e+00 1.12357063e-02-3.13558070e-06 1.59502818e-10 3.01357560e-14    2
-5.57414981e+04-1.53809923e+01 3.13168541e-01 3.25739975e-02-2.58358905e-05    3
 1.08925098e-08-1.87287967e-12-5.36203653e+04 2.34914872e+01                   4
CH3NO                   C   1H   3O   1N   1G    300.00   3500.00  860.00      1
 1.73828229e+00 1.65479495e-02-8.69271695e-06 2.17002760e-09-2.08463444e-13    2
 8.36473513e+03 1.74966005e+01 2.23451684e+00 1.42398818e-02-4.66701756e-06    3
-9.50669597e-10 6.98715974e-13 8.27938279e+03 1.51773992e+01                   4
CH3NO2                  C   1H   3O   2N   1G    300.00   3500.00 1620.00      1
 5.94771391e+00 1.22319078e-02-4.98716389e-06 9.73177561e-10-7.54873508e-14    2
-1.14691242e+04-2.73415041e+00-2.05952276e-01 2.74261453e-02-1.90559023e-05    3
 6.76278185e-09-9.68944802e-13-9.47533640e+03 2.99224212e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00  700.00      1
 6.88420582e-01 1.44971301e-02-7.59068052e-06 1.92522389e-09-1.90011116e-13    2
 1.18330404e+03 1.95838279e+01 2.13962537e+00 6.20453130e-03 1.01791740e-05    3
-1.49984471e-08 5.85415708e-12 9.80135371e+02 1.31002120e+01                   4
CH3OCH2                 C   2H   5O   1     G    300.00   3500.00  750.00      1
 2.76373432e+00 2.09427776e-02-1.03906311e-05 2.45853855e-09-2.25935821e-13    2
-6.59718889e+02 1.23154396e+01 2.98724171e+00 1.97507382e-02-8.00655224e-06    3
 3.39357381e-10 4.80457902e-13-6.93244997e+02 1.13014447e+01                   4
CH3OCH3                 C   2H   6O   1     G    300.00   3500.00  700.00      1
 8.15389478e-01 2.72675400e-02-1.40181429e-05 3.43685384e-09-3.25542356e-13    2
-2.31745898e+04 1.99239256e+01 1.74097325e+00 2.19784899e-02-2.68446400e-06    3
-7.35712603e-09 3.52945045e-12-2.33041715e+04 1.57886515e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 2.14769740e+00 2.46740524e-02-1.35238094e-05 3.44782067e-09-3.34980467e-13    2
-4.40372636e+04 1.69024645e+01 3.51192337e+00 1.68784755e-02 3.18099831e-06    3
-1.24615200e-08 5.34692693e-12-4.42282552e+04 1.08074480e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849390e-09-3.11411020e-13    2
-2.07085510e+04 1.59117693e+01 4.66126893e+00 9.68655554e-03 1.14715528e-05    3
-1.83003965e-08 7.03409939e-12-2.10131064e+04 6.50453092e+00                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00  700.00      1
 9.34193000e-01 1.60266556e-02-8.00101466e-06 1.97129714e-09-1.91599484e-13    2
-2.50979789e+04 1.91008457e+01 2.88895785e+00 4.85657077e-03 1.59348814e-05    3
-2.08247943e-08 7.94986176e-12-2.53716460e+04 1.03674509e+01                   4
CH3ONO                  C   1H   3O   2N   1G    300.00   3500.00 1800.00      1
 8.58034518e+00 8.90954082e-03-3.35922089e-06 6.18588139e-10-4.68096982e-14    2
-1.15569624e+04-1.97194056e+01 1.99249583e+00 2.35492060e-02-1.55589419e-05    3
 5.13700333e-09-6.74367363e-13-9.18533663e+03 1.59354094e+01                   4
CH3ONO2                 C   1H   3O   3N   1G    300.00   3500.00 1800.00      1
 1.07457798e+01 1.03362024e-02-4.39539782e-06 8.95959797e-10-7.26862027e-14    2
-1.81031090e+04-3.08875015e+01 1.35155390e+00 3.12122600e-02-2.17921125e-05    3
 7.33918744e-09-9.67578931e-13-1.47211877e+04 1.99560088e+01                   4
CH3OO                   C   1H   3O   2     G    300.00   3500.00 1300.00      1
 3.46521970e+00 1.23938518e-02-5.59614682e-06 1.22616716e-09-1.06238815e-13    2
 6.86982281e+02 1.04298931e+01 4.30117244e+00 9.82168948e-03-2.62826727e-06    3
-2.95822349e-10 1.86451475e-13 4.69634569e+02 6.17758023e+00                   4
CH3OOH                  C   1H   4O   2     G    300.00   3500.00 1800.00      1
 5.50146514e+00 1.13975421e-02-3.82130848e-06 4.38704910e-10-2.90617476e-15    2
-1.79784234e+04-4.65581411e-01 5.93430876e+00 1.04356674e-02-3.01974623e-06    3
 1.41830001e-10 3.83264515e-14-1.81342471e+04-2.80822136e+00                   4
CH4                     C   1H   4          G    300.00   3500.00 1070.00      1
-2.82321416e-01 1.42739336e-02-6.77628877e-06 1.55380951e-09-1.39473841e-13    2
-9.36383584e+03 2.03507024e+01 2.85765313e+00 2.53571100e-03 9.67916346e-06    3
-8.69880870e-09 2.25599770e-12-1.00357904e+04 4.98969392e+00                   4
CHCHCH3                 C   3H   5          G    300.00   3500.00 1800.00      1
 1.00124373e+01 7.55815802e-03-1.17096962e-06-2.01794819e-10 4.72987983e-14    2
 2.78641947e+04-2.75169832e+01 6.10512020e-01 2.84513252e-02-1.85819423e-05    3
 6.24671358e-09-8.48327368e-13 3.12488878e+04 2.33681976e+01                   4
CN                      C   1N   1          G    300.00   3500.00  810.00      1
 2.73859606e+00 2.23580966e-03-1.33797023e-06 4.34996429e-10-5.05222621e-14    2
 5.14568835e+04 8.20480076e+00 4.08532688e+00-4.41471288e-03 1.09778123e-05    3
-9.70145006e-09 3.07801060e-12 5.12387131e+04 1.99138758e+00                   4
CO                      C   1O   1          G    300.00   3500.00 1000.00      1
 2.68595014e+00 2.12486373e-03-1.04548608e-06 2.45538864e-10-2.22550981e-14    2
-1.41423615e+04 7.96579426e+00 3.81890943e+00-2.40697343e-03 5.75226966e-06    3
-4.28629830e-09 1.11070419e-12-1.43689533e+04 2.49992060e+00                   4
CO2                     C   1O   2          G    300.00   3500.00 1620.00      1
 5.07830985e+00 2.05366041e-03-5.94311265e-07 5.38675131e-11 1.66346855e-15    2
-4.92442103e+04-4.47815290e+00 2.44892797e+00 8.54596135e-03-6.60570102e-06    3
 2.52769046e-09-3.80099332e-13-4.83922906e+04 9.47557732e+00                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155283e-02-1.38949871e-05 2.56768166e-09-1.71519559e-13    2
-2.17187243e+04-3.95715124e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733025e-12-1.73470426e+04 4.54334869e+01                   4
CSOLID                  C   1               G    300.00   3500.00 1470.00      1
 1.73007911e+00 1.24133836e-03-3.99676695e-07 5.50148663e-11-1.79078883e-15    2
-8.17038240e+02-1.00735633e+01-8.82758554e-01 8.35110072e-03-7.65453624e-06    3
 3.34520060e-09-5.61346186e-13-4.88639663e+01 3.53849619e+00                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459579e+00 2.39841575e-02-8.32755388e-06 8.47127653e-10 2.86249484e-14    2
 3.08659308e+03-9.73181554e+00-5.14379339e+00 6.04552342e-02-5.17455024e-05    3
 2.38195872e-08-4.52940274e-12 5.98166715e+03 4.83481227e+01                   4
CYC5H5                  C   5H   5          G    300.00   3500.00  700.00      1
 4.01652575e+00 2.68451891e-02-1.26423018e-05 2.78092332e-09-2.35299436e-13    2
 2.91110159e+04 1.44025794e+00-2.58737408e+00 6.45817595e-02-9.35063814e-05    3
 7.97943325e-08-2.77400884e-11 3.00355619e+04 3.09448116e+01                   4
CYC5H6                  C   5H   6          G    300.00   3500.00 1020.00      1
 1.70141558e+00 3.79065957e-02-2.19495256e-05 6.12706526e-09-6.63672518e-13    2
 1.38484401e+04 1.22453451e+01-6.32922867e+00 6.93993183e-02-6.82623529e-05    3
 3.63968870e-08-8.08274648e-12 1.54866915e+04 5.11475893e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099915e+00 2.71082714e-02-1.07932862e-05 1.95387666e-09-1.31111174e-13    2
-1.09862538e+03-2.37608447e+01-6.56863980e+00 6.82031726e-02-5.30140751e-05    3
 2.12327757e-08-3.43229252e-12 3.28126920e+03 5.42801525e+01                   4
CYC6-OO                 C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.87814621e+01 3.54361927e-02-1.49718784e-05 3.04328287e-09-2.46478319e-13    2
-1.95252830e+04-7.87240875e+01-6.50623568e+00 9.16310766e-02-6.18009483e-05    3
 2.03873828e-08-2.65538109e-12-1.04217118e+04 5.81382079e+01                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283791e-14    2
-3.55499047e+04-1.30447295e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.49648189e+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.17655243e+01 3.67451404e-02-1.42717448e-05 2.74140449e-09-2.13135508e-13    2
-3.59903393e+04-5.10812501e+01-1.06696444e+01 9.82113560e-02-7.74219664e-05    3
 3.15771221e-08-5.15075839e-12-2.94392700e+04 6.56457555e+01                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.91587814e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.29538877e+01                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.91384147e+01 3.64873063e-02-1.63612962e-05 3.53264562e-09-3.02111689e-13    2
-1.43294351e+04-7.86383640e+01-4.87015408e+00 8.98396814e-02-6.08216088e-05    3
 1.99994281e-08-2.58916481e-12-5.68635037e+03 5.13010187e+01                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624858e+01 2.76360017e-02-1.05259858e-05 1.89586361e-09-1.35054773e-13    2
-9.29985245e+03-6.25064559e+01-6.01517655e+00 7.46974737e-02-4.97438791e-05    3
 1.64210093e-08-2.15243611e-12-1.67589399e+03 5.21114707e+01                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.29323176e+01 2.20056554e-02-7.35242348e-06 1.07816406e-09-5.64635915e-14    2
-2.79806200e+04-1.10525204e+02-1.05629257e+01 9.64395294e-02-6.93806518e-05    3
 2.40515820e-08-3.24721608e-12-1.59223324e+04 7.07580407e+01                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.18028612e+01 2.41377428e-02-8.73118284e-06 1.46035609e-09-9.51866870e-14    2
-2.87387454e+04-1.06217525e+02-1.25990095e+01 1.00586344e-01-7.24383509e-05    3
 2.50556035e-08-3.37230438e-12-1.63540719e+04 7.99725758e+01                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.14079592e+01 2.50825461e-02-9.38039634e-06 1.64525432e-09-1.14247640e-13    2
-3.89741817e+04-1.05728233e+02-1.45960517e+01 1.05091459e-01-7.60544907e-05    3
 2.63393633e-08-3.54398500e-12-2.60127378e+04 8.91329846e+01                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.15965428e+01 4.02887933e-02-1.86685839e-05 4.15568433e-09-3.64030709e-13    2
-3.62221493e+04-4.27468434e+01-6.46490379e+00 8.04253413e-02-5.21157073e-05    3
 1.65435078e-08-2.08456175e-12-2.97200285e+04 5.50054734e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879190e+01 3.94798364e-02-1.80474738e-05 3.97976998e-09-3.47933573e-13    2
 4.69934406e+02-4.15743644e+01-9.20200373e+00 8.50129981e-02-5.59917752e-05    3
 1.80332150e-08-2.29980093e-12 7.84630661e+03 6.93213721e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578097e+01 4.34354098e-02-2.02455774e-05 4.54245292e-09-4.01195170e-13    2
-2.30439963e+04-4.47863376e+01-9.43363126e+00 8.94163897e-02-5.85630607e-05    3
 1.87341134e-08-2.37225913e-12-1.55950776e+04 6.72000574e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772260e+00 3.45074855e-02-1.63846780e-05 3.69260975e-09-3.24421026e-13    2
 5.74022139e+03-2.73566208e+01-6.91358136e+00 7.63364895e-02-5.84944135e-05    3
 2.25336547e-08-3.48567018e-12 1.03834500e+04 5.40276160e+01                   4
CYC6H9                  C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670463e+01 2.75651338e-02-1.13337615e-05 2.23021652e-09-1.74683445e-13    2
 7.93866332e+03-5.85441979e+01-6.48639356e+00 7.34616669e-02-4.95808724e-05    3
 1.63958131e-08-2.14212742e-12 1.53739017e+04 5.32365273e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525256e+01 3.24730728e-02-1.15459374e-05 1.79679054e-09-9.97833662e-14    2
-5.30753651e+03-1.13355893e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932248e-08-9.37220078e-12 5.02765510e+03 7.60497478e+01                   4
DIFENET                 C  12H  10O   1     G    300.00   3500.00 1430.00      1
 1.71548107e+01 5.25374196e-02-2.45657222e-05 5.58244776e-09-4.99409896e-13    2
-3.29704394e+03-6.49985669e+01-8.57458099e+00 1.24507746e-01-1.00059071e-04    3
 4.07774824e-08-6.65238798e-12 4.06156207e+03 6.83336207e+01                   4
DIPE                    C   6H  14O   1     G    300.00   3500.00 1380.00      1
 1.11573928e+01 4.99175659e-02-2.25561386e-05 4.38444843e-09-3.06549364e-13    2
-4.59357929e+04-3.06117763e+01-2.50745274e+00 8.95258138e-02-6.56085820e-05    3
 2.51827303e-08-4.07435404e-12-4.21642955e+04 3.97144256e+01                   4
DME-OO                  C   2H   5O   3     G    300.00   3500.00  870.00      1
 3.58974575e+00 2.80960123e-02-1.49224205e-05 3.71355557e-09-3.53703711e-13    2
-1.93352293e+04 1.47278303e+01 5.41345468e+00 1.97111437e-02-4.65750394e-07    3
-7.36435253e-09 2.82960321e-12-1.96525546e+04 6.18346241e+00                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   3500.00 1800.00      1
 9.57989146e+00 2.53360331e-02-1.13706887e-05 2.45690684e-09-2.09295699e-13    2
-3.48199648e+04-1.16031904e+01 7.85487749e+00 2.91693975e-02-1.45651591e-05    3
 3.64004400e-09-3.73620304e-13-3.41989598e+04-2.26705495e+00                   4
DME-OQOOH               C   2H   4O   4     G    300.00   3500.00 1760.00      1
 1.54960865e+01 1.58758106e-03 2.24425901e-06-9.74237206e-10 1.03773065e-13    2
-4.69655432e+04-5.18401164e+01 3.62388957e+00 2.85698467e-02-2.07519902e-05    3
 7.73646324e-09-1.13354234e-12-4.27865299e+04 1.21478877e+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   3500.00 1800.00      1
 9.52551493e+00 1.89562856e-02-9.27557330e-06 2.15192754e-09-1.93905680e-13    2
-1.72537528e+04-1.74698518e+01 5.12252607e+00 2.87407053e-02-1.74292564e-05    3
 5.17181016e-09-6.13333823e-13-1.56686768e+04 6.36004246e+00                   4
DMF                     C   6H   8O   1     G    300.00   3500.00 1590.00      1
 1.38889506e+01 2.49736923e-02-8.98421021e-06 1.42738238e-09-7.97717945e-14    2
-2.20872034e+04-4.94041109e+01-2.31533181e+00 6.57391826e-02-4.74422199e-05    3
 1.75523340e-08-2.61514155e-12-1.69342416e+04 3.62866615e+01                   4
DMF-3YL                 C   6H   7O   1     G    300.00   3500.00 1620.00      1
 1.41703395e+01 2.18230092e-02-7.69511407e-06 1.17891300e-09-6.12376638e-14    2
 1.19557792e+04-4.86583489e+01-1.12307984e+00 5.95845385e-02-4.26594930e-05    3
 1.55675463e-08-2.28170577e-12 1.69108471e+04 3.25015043e+01                   4
ERC4H8CHO               C   5H   9O   1     G    300.00   3500.00  750.00      1
-3.04813054e-01 5.67977502e-02-3.24057642e-05 8.50471985e-09-8.41763290e-13    2
-5.21420511e+03 3.41933259e+01 6.22525332e+00 2.19707295e-02 3.72482771e-05    3
-5.34099835e-08 1.97964712e-11-6.19371507e+03 4.56811339e+00                   4
ETBE                    C   6H  14O   1     G    300.00   3500.00 1280.00      1
 1.16559136e+01 4.67933987e-02-1.93342014e-05 3.59185140e-09-2.45564975e-13    2
-4.60322114e+04-3.38084939e+01-3.48005604e+00 9.40933039e-02-7.47637778e-05    3
 3.24614225e-08-5.88415307e-12-4.21574031e+04 4.29502770e+01                   4
ETC3H4O2                C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920429e+01 1.38871300e-02-6.12561993e-06 1.30548845e-09-1.09965765e-13    2
-3.57026988e+04-2.69350036e+01 1.17378045e-01 4.67086294e-02-4.58290467e-05    3
 2.26514168e-08-4.41358036e-12-3.31793820e+04 2.43405589e+01                   4
ETEROMD                 C  11H  20O   3     G    300.00   3500.00 1760.00      1
 4.14249213e+01 4.51122053e-02-1.56530088e-05 2.49214075e-09-1.50324737e-13    2
-8.95581279e+04-1.84296546e+02-1.24327962e-01 1.39542317e-01-9.61332178e-05    3
 3.29770684e-08-4.48057014e-12-7.49327921e+04 3.96429285e+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   3500.00 1310.00      1
 4.32126695e+01 9.17256499e-02-3.02788098e-05 4.53882493e-09-2.50045022e-13    2
-1.06117741e+05-1.75617618e+02-8.73011664e+00 2.50329577e-01-2.11886360e-04    3
 9.69599701e-08-1.78876681e-11-9.25087311e+04 8.90022613e+01                   4
ETMB583                 C   5H   8O   3     G    300.00   3500.00 1270.00      1
 1.75630365e+01 2.35383857e-02-7.56913166e-06 1.05837457e-09-4.95698273e-14    2
-6.27369638e+04-6.15054259e+01-4.60165685e+00 9.33484435e-02-9.00219559e-05    3
 4.43406970e-08-8.56971204e-12-5.71071317e+04 5.07241435e+01                   4
FLUORENE                C  13H  10          G    300.00   3500.00 1440.00      1
 2.91248872e+01 2.85362024e-02-5.66199729e-06-5.67026725e-10 1.91134972e-13    2
 9.75119358e+03-1.37159218e+02-1.43465120e+01 1.49290089e-01-1.31447296e-04    3
 5.76669078e-08-9.91892310e-12 2.22709565e+04 8.84167006e+01                   4
GLIET                   C   2H   6O   2     G    300.00   3500.00 1470.00      1
 6.66621468e+00 1.87459315e-02-7.66039208e-06 1.53874843e-09-1.24203245e-13    2
-4.95959120e+04-6.01671900e+00 9.46220545e-01 3.43105414e-02-2.35426471e-05    3
 8.74158516e-09-1.34917548e-12-4.79142337e+04 2.37826449e+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   3500.00 1290.00      1
 1.14796489e+01 2.36292461e-02-8.98384419e-06 1.70355137e-09-1.31527258e-13    2
-7.41781076e+04-2.56707288e+01 1.97850806e-01 5.86115658e-02-4.96609601e-05    3
 2.27253167e-08-4.20551279e-12-7.12674037e+04 3.16302477e+01                   4
H                       H   1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
 2.54716200e+04-4.60117600e-01 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25 2.54716200e+04-4.60117600e-01                   4
H2                      H   2               G    300.00   3500.00  750.00      1
 3.73110902e+00-8.86706214e-04 1.12286897e-06-3.74349782e-10 4.17963674e-14    2
-1.08851547e+03-5.35285855e+00 3.08866003e+00 2.53968841e-03-5.72992027e-06    3
 5.71701843e-09-1.98865970e-12-9.92148124e+02-2.43823459e+00                   4
H2CN                    C   1H   2N   1     G    300.00   3500.00 1800.00      1
 5.22111320e+00 3.42647499e-03-8.36137799e-07 4.74833030e-11 4.28153350e-15    2
 2.75312364e+04-4.80262216e+00 1.81354567e+00 1.09988473e-02-7.14644805e-06    3
 2.38463525e-09-3.20322903e-13 2.87579607e+04 1.36398442e+01                   4
H2NO                    H   2O   1N   1     G    300.00   3500.00 1200.00      1
 1.43405821e+00 9.01333883e-03-3.38828321e-06 4.28655869e-10-2.36936075e-15    2
 7.27341661e+03 1.79341864e+01 2.78935895e+00 4.49566971e-03 2.25880318e-06    3
-2.70861435e-09 6.51228601e-13 6.94814443e+03 1.11485432e+01                   4
H2O                     H   2O   1          G    300.00   3500.00 1590.00      1
 2.30940463e+00 3.65433887e-03-1.22983871e-06 2.11931683e-10-1.50333493e-14    2
-2.97294901e+04 8.92765177e+00 4.03530937e+00-6.87559833e-04 2.86629214e-06    3
-1.50552360e-09 2.55006790e-13-3.02783278e+04-1.99201641e-01                   4
H2O2                    H   2O   2          G    300.00   3500.00 1180.00      1
 4.56163072e+00 4.35560969e-03-1.48694629e-06 2.38275424e-10-1.46610352e-14    2
-1.80016693e+04 5.66597119e-01 2.91896355e+00 9.92397296e-03-8.56537418e-06    3
 4.23738723e-09-8.61930485e-13-1.76139998e+04 8.76340177e+00                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1800.00      1
 7.44900312e+00 1.01177830e-03 3.02918165e-07-2.13909391e-10 2.81815208e-14    2
 1.86458955e+04-1.30987733e+01 4.44514163e+00 7.68702606e-03-5.25978830e-06    3
 1.84635226e-09-2.57965931e-13 1.97272856e+04 3.15875175e+00                   4
HCN                     C   1H   1N   1     G    300.00   3500.00  850.00      1
 3.48152100e+00 3.81748410e-03-1.53642929e-06 3.02291150e-10-2.35861473e-14    2
 1.50427831e+04 3.30702298e+00 2.53139665e+00 8.28865751e-03-9.42673531e-06    3
 6.49076646e-09-1.84372594e-12 1.52043042e+04 7.73641055e+00                   4
HCNO                    C   1H   1O   1N   1G    300.00   3500.00 1350.00      1
 7.12423974e+00 1.61853378e-03 2.31339437e-07-2.53211924e-10 3.63453797e-14    2
 1.67567928e+04-1.48886865e+01 2.20954024e+00 1.61806064e-02-1.59487412e-05    3
 7.73695136e-09-1.44331449e-12 1.80837616e+04 1.02968215e+01                   4
HCO                     C   1H   1O   1     G    300.00   3500.00  920.00      1
 2.44772078e+00 5.65570555e-03-3.01329556e-06 7.57702524e-10-7.26129631e-14    2
 4.31149160e+03 1.15871953e+01 3.74218864e+00 2.75844059e-05 6.16298892e-06    3
-5.89177898e-09 1.73431136e-12 4.07330951e+03 5.45007090e+00                   4
HCO3                    C   1H   1O   3     G    300.00   3500.00 1800.00      1
 5.04067718e+00 8.66656109e-03-4.28958277e-06 1.00563376e-09-9.13599886e-14    2
-1.77902136e+04 5.78191516e+00 3.79300672e+00 1.14391621e-02-6.60008362e-06    3
 1.86137482e-09-2.10212913e-13-1.73410522e+04 1.25345680e+01                   4
HCO3H                   C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230668e+01 4.43563253e-03-1.56188514e-06 2.43424395e-10-1.38391379e-14    2
-3.81313332e+04-2.33590722e+01 2.47434199e+00 2.16898607e-02-1.63512235e-05    3
 5.87745807e-09-8.18701091e-13-3.54892796e+04 1.72835470e+01                   4
HCOOH                   C   1H   2O   2     G    300.00   3500.00 1800.00      1
 5.80573302e+00 6.82017393e-03-2.95480608e-06 6.14340060e-10-5.06753135e-14    2
-4.80534416e+04-6.42993389e+00 1.36256505e+00 1.66938805e-02-1.11828949e-05    3
 3.66178037e-09-4.73930912e-13-4.64539011e+04 1.76174180e+01                   4
HE                      HE  1               G    300.00   3500.00 1490.00      1
 2.50000000e+00 7.40336223e-15-5.56967416e-18 1.73924876e-21-1.92673709e-25    2
-7.45375000e+02 9.28723974e-01 2.50000000e+00-4.07455160e-15 5.98527266e-18    3
-3.43074982e-21 6.74775716e-25-7.45375000e+02 9.28723974e-01                   4
HNCO                    C   1H   1O   1N   1G    300.00   3500.00 1660.00      1
 7.29502452e+00 4.88032844e-04 8.74568316e-07-4.09105701e-10 5.01959355e-14    2
-1.52722297e+04-1.41696888e+01 2.99127956e+00 1.08585026e-02-8.49633812e-06    3
 3.35431054e-09-5.16583618e-13-1.38433864e+04 8.77460657e+00                   4
HNNO                    H   1O   1N   2     G    300.00   3500.00 1360.00      1
 4.88500308e+00 5.60936901e-03-2.60717829e-06 5.93839036e-10-5.41495114e-14    2
 2.58926738e+04 6.01980007e-01 2.29344827e+00 1.32315890e-02-1.10140386e-05    3
 4.71484900e-09-8.11688108e-13 2.65975767e+04 1.39015974e+01                   4
HNO                     H   1O   1N   1     G    300.00   3500.00  900.00      1
 2.72673666e+00 5.06770488e-03-2.61122761e-06 6.38493559e-10-6.01581004e-14    2
 1.09769405e+04 9.63912842e+00 3.40204752e+00 2.06632330e-03 2.39107502e-06    3
-3.06691580e-09 9.69122277e-13 1.08553846e+04 6.45229501e+00                   4
HNO2                    H   1O   2N   1     G    300.00   3500.00 1800.00      1
 3.30359406e+00 7.74006618e-03-3.91474332e-06 9.47112178e-10-8.88494507e-14    2
-8.65702544e+03 7.10072496e+00 1.68890715e+00 1.13282593e-02-6.90490427e-06    3
 2.05457920e-09-2.42664314e-13-8.07573815e+03 1.58397474e+01                   4
HO2                     H   1O   2          G    300.00   3500.00 1540.00      1
 4.16318067e+00 1.99798265e-03-4.89192086e-07 7.71153172e-11-7.30772104e-15    2
 4.41348948e+01 2.95517985e+00 2.85241381e+00 5.40257188e-03-3.80535043e-06    3
 1.51268170e-09-2.40354212e-13 4.47851086e+02 9.84483831e+00                   4
HOCN                    C   1H   1O   1N   1G    300.00   3500.00 1760.00      1
 6.92286755e+00 1.77083687e-04 1.06417841e-06-4.55819441e-10 5.43563991e-14    2
-3.77375638e+03-1.08544042e+01 3.05788784e+00 8.96112848e-03-6.42222341e-06    3
 2.37993882e-09-3.48450172e-13-2.41328352e+03 9.97681509e+00                   4
HONO                    H   1O   2N   1     G    300.00   3500.00 1420.00      1
 5.88742112e+00 3.49329101e-03-1.17730803e-06 1.65569378e-10-6.87715202e-15    2
-1.14386309e+04-5.23866548e+00 2.37883184e+00 1.33766411e-02-1.16174666e-05    3
 5.06705227e-09-8.69814280e-13-1.04421916e+04 1.29185606e+01                   4
HONO2                   H   1O   3N   1     G    300.00   3500.00 1310.00      1
 5.20949091e+00 9.97123440e-03-5.50725421e-06 1.39250696e-09-1.33157469e-13    2
-1.74464288e+04-1.35430787e+00 8.85706040e-01 2.31736309e-02-2.06245022e-05    3
 9.08576291e-09-1.60133609e-12-1.63135971e+04 2.06729940e+01                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1420.00      1
 4.21122112e+01 1.11834123e-01-5.11978482e-05 1.12541459e-08-9.72533984e-13    2
-7.89343498e+04-1.80495570e+02-6.54289827e+00 2.48890769e-01-1.95975996e-04    3
 7.92251073e-08-1.29392525e-11-6.51162987e+04 7.12984570e+01                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1590.00      1
 5.03105902e+01 8.85535013e-02-3.63077668e-05 7.13747183e-09-5.56692148e-13    2
-1.01978074e+05-2.30341253e+02-5.93668664e+00 2.30056085e-01-1.69800770e-04    3
 6.31093809e-08-9.35730677e-12-8.40914402e+04 6.71031189e+01                   4
IC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1460.00      1
 4.22439745e+01 1.02589738e-01-4.54459633e-05 9.70909447e-09-8.19911243e-13    2
-6.26654622e+04-1.86283114e+02-7.79323360e+00 2.39677979e-01-1.86290047e-04    3
 7.40214614e-08-1.18323028e-11-4.80545975e+04 7.40533932e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453588e+01 7.53296743e-02-2.79263242e-05 4.92908201e-09-3.44364401e-13    2
-5.61938874e+04-2.43048234e+02-8.95216175e+00 2.21020633e-01-1.60372651e-04    3
 5.84427492e-08-8.45249579e-12-3.63617056e+04 7.69829165e+01                   4
IC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1460.00      1
 3.94749769e+01 1.06211481e-01-4.74108472e-05 1.02029370e-08-8.67107397e-13    2
-6.81954459e+04-1.73182708e+02-7.55515778e+00 2.35061165e-01-1.79790660e-04    3
 7.06503399e-08-1.12176901e-11-5.44626465e+04 7.15084222e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524600e+01 8.54680758e-02-3.36612723e-05 6.38202029e-09-4.82094887e-13    2
-7.78744143e+04-2.24182950e+02-9.93612250e+00 2.29338723e-01-1.69388298e-04    3
 6.32906266e-08-9.42998897e-12-5.96884450e+04 7.82391931e+01                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   3500.00 1370.00      1
 4.07769110e+01 1.15135971e-01-5.36319133e-05 1.19826916e-08-1.04989886e-12    2
-8.16821240e+04-1.74509322e+02-7.08781179e+00 2.54886986e-01-2.06643974e-04    3
 8.64411154e-08-1.46372025e-11-6.85671899e+04 7.14786263e+01                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   3500.00 1560.00      1
 5.03537527e+01 8.72534729e-02-3.55849544e-05 6.99643634e-09-5.47405935e-13    2
-6.86134004e+04-2.32227161e+02-7.33743336e+00 2.35179591e-01-1.77821606e-04    3
 6.77813303e-08-1.02885748e-11-5.06137504e+04 7.17539151e+01                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1220.00      1
 1.23035624e+01 2.79964883e-02-1.33482910e-05 3.03524083e-09-2.69271163e-13    2
-2.25784829e+04-2.78550798e+01 1.73143843e+00 6.26591900e-02-5.59663668e-05    3
 2.63238068e-08-5.04151829e-12-1.99988847e+04 2.52515831e+01                   4
IC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1270.00      1
 1.04498043e+01 2.29490980e-02-1.05757759e-05 2.34172678e-09-2.03669153e-13    2
-5.22299426e+03-2.40008692e+01-1.71110880e-01 5.64007993e-02-5.00856593e-05    3
 2.30818231e-08-4.28636527e-12-2.52528181e+03 2.97774852e+01                   4
IC3H5CHO                C   4H   6O   1     G    300.00   3500.00 1370.00      1
 8.96605760e+00 2.20962385e-02-1.00901145e-05 2.22139279e-09-1.91792264e-13    2
-1.79920102e+04-2.11939239e+01 6.92941977e-01 4.62513206e-02-3.65372847e-05    3
 1.50910620e-08-2.54027204e-12-1.57251765e+04 2.13235423e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1630.00      1
 8.48779790e+00 1.53259253e-02-4.76474417e-06 3.92065263e-10 2.47111520e-14    2
 5.50507422e+03-2.12719618e+01 2.73725246e-01 3.54831588e-02-2.33143455e-05    3
 7.97881429e-09-1.13890066e-12 8.18286190e+03 2.23694223e+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.25375038e+01 2.06759832e-02-7.90606663e-06 1.44761601e-09-1.05776578e-13    2
-3.22363635e+04-4.10505202e+01-3.44732114e-01 4.93031741e-02-3.17620591e-05    3
 1.02831688e-08-1.33293668e-12-2.75987585e+04 2.86708279e+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1310.00      1
 6.28069615e+00 2.59370043e-02-1.05350747e-05 1.92921360e-09-1.30183993e-13    2
-3.63768639e+04-6.66341882e+00-3.00574060e-01 4.60324859e-02-3.35451681e-05    3
 1.36391848e-08-2.36491132e-12-3.46525711e+04 2.68645272e+01                   4
IC3H7OO                 C   3H   7O   2     G    300.00   3500.00 1260.00      1
 7.34738699e+00 2.68252330e-02-1.24179691e-05 2.76645854e-09-2.42147350e-13    2
-1.06484855e+04-8.92587196e+00 1.07341266e+00 4.67426118e-02-3.61291344e-05    3
 1.53120486e-08-2.73135173e-12-9.06744395e+03 2.27924165e+01                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1570.00      1
 1.51567879e+01 2.57227734e-02-1.11020451e-05 2.28943519e-09-1.86269530e-13    2
-4.30658407e+04-4.59845002e+01 9.69279340e-01 6.18692920e-02-4.56369355e-05    3
 1.69539322e-08-2.52138051e-12-3.86109630e+04 2.88616666e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955794e+00 3.23747266e-02-1.18655436e-05 1.37455178e-09 1.57073476e-14    2
-1.97025810e+04-6.34483422e+00-1.85965328e+00 5.58007940e-02-3.97537190e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177121e+00 3.67769036e-02-1.77031336e-05 3.74786262e-09-2.92191280e-13    2
 1.31214242e+04 2.00120538e+01 3.86129991e+00 2.14653110e-02 1.51074220e-05    3
-2.75002856e-08 1.08678616e-11 1.27462902e+04 8.04059744e+00                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385768e+03-1.72949366e+01 7.17301598e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035734e-13-3.72372397e+03 2.01415164e+01                   4
IC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.44537517e+01 2.20810695e-02-7.57959310e-06 1.19533670e-09-7.16167606e-14    2
-4.15822810e+04-5.13315495e+01-5.45479447e-01 5.54126942e-02-3.53559470e-05    3
 1.14828752e-08-1.50044155e-12-3.61825578e+04 2.98474183e+01                   4
IC4H9P                  C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221491e-06 8.09648923e-10 4.02033219e-14    2
 3.37759298e+03-1.61084037e+01-1.15582376e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   3500.00 1380.00      1
 8.54295826e+00 3.45220773e-02-1.59311943e-05 3.53852672e-09-3.08950056e-13    2
-1.29532173e+04-1.39825068e+01 7.00555201e-01 5.72536803e-02-4.06394585e-05    3
 1.54748862e-08-2.47133403e-12-1.07887140e+04 2.63784632e+01                   4
IC4H9T                  C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871688e+00 2.55264450e-02-8.65284050e-06 8.24419704e-10 3.80550653e-14    2
 8.35470581e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397360e-05    3
 1.42467509e-08-2.35878979e-12 3.41363196e+03 3.01901373e+01                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   3500.00 1260.00      1
 9.11667611e+00 3.41757258e-02-1.58797345e-05 3.54686464e-09-3.10976548e-13    2
-1.64591648e+04-1.96564028e+01 4.84069009e-01 6.15808277e-02-4.85048558e-05    3
 2.08088336e-08-3.73597039e-12-1.42837478e+04 2.39860330e+01                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1290.00      1
 1.30518446e+01 3.65484801e-02-1.74274782e-05 3.96741952e-09-3.52552034e-13    2
-2.47096139e+04-3.04334702e+01 1.64511788e+00 7.19181753e-02-5.85550308e-05    3
 2.52219686e-08-4.47165070e-12-2.17666784e+04 2.75020267e+01                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   3500.00 1350.00      1
 1.14809469e+01 3.08095616e-02-1.41939360e-05 3.14755455e-09-2.74422165e-13    2
-7.45268236e+03-2.80879239e+01-1.93281563e-01 6.53998681e-02-5.26276099e-05    3
 2.21271466e-08-3.78916143e-12-4.30064068e+03 3.17369695e+01                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1240.00      1
 1.39939782e+01 3.54845222e-02-1.68915059e-05 3.83671077e-09-3.40131614e-13    2
-2.83614519e+04-3.70531088e+01 1.55094393e+00 7.56233424e-02-6.54465303e-05    3
 2.99415626e-08-5.60320657e-12-2.52755794e+04 2.56539769e+01                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   3500.00 1270.00      1
 1.20890742e+01 3.03954175e-02-1.40883982e-05 3.13822121e-09-2.74437748e-13    2
-1.09705556e+04-3.28537329e+01-4.26302143e-01 6.98139255e-02-6.06456912e-05    3
 2.75777451e-08-5.08536764e-12-7.79165002e+03 3.05171096e+01                   4
IC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 2.13459841e+01 8.88367161e-03 1.59648418e-06-1.31808203e-09 1.74600856e-13    2
-1.26620076e+04-8.94699897e+01-1.59634535e+00 5.98666259e-02-4.08893110e-05    3
 1.44173977e-08-2.01088244e-12-4.40276906e+03 3.46986831e+01                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   3500.00 1710.00      1
 3.48314225e+01 3.98146097e-02-1.43978345e-05 2.42273589e-09-1.57988116e-13    2
-5.01227380e+04-1.45334518e+02 1.76391327e+00 1.17165508e-01-8.22495000e-05    3
 2.88756269e-08-4.02536985e-12-3.88136498e+04 3.19375985e+01                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   3500.00 1770.00      1
 3.33140926e+01 3.48304479e-02-1.19632189e-05 1.85711682e-09-1.07309433e-13    2
-6.88276671e+04-1.40834098e+02 5.55148980e-01 1.08861959e-01-7.47017874e-05    3
 2.54874628e-08-3.44492892e-12-5.72310011e+04 3.59135548e+01                   4
IC8-QOOH                C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574275e-02-1.91478836e-05 3.78861311e-09-2.97862012e-13    2
-2.91331926e+04-1.00455337e+02-9.92411236e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616063e+01 4.14292819e-02-1.28170544e-05 1.66806736e-09-6.58961711e-14    2
-2.24684067e+04-7.38514296e+01-5.35586581e+00 1.10622059e-01-8.69521729e-05    3
 3.69705048e-08-6.36990285e-12-1.56875145e+04 5.11323811e+01                   4
IC8H16O                 C   8H  16O   1     G    300.00   3500.00 1730.00      1
 2.92525449e+01 3.42835226e-02-1.16024061e-05 1.77291874e-09-1.00401812e-13    2
-4.92824114e+04-1.33818841e+02-8.05235857e+00 1.20537635e-01-8.63892084e-05    3
 3.05924957e-08-4.26508057e-12-3.63749148e+04 6.66033697e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104230e+01 3.01796816e-02-5.82184991e-06 1.42085860e-11 7.60110759e-14    2
-1.80373025e+04-1.14981197e+02-3.32961207e+00 1.08192845e-01-8.23053435e-05    3
 3.33403496e-08-5.36943680e-12-8.90625182e+03 4.16697269e+01                   4
IC8H17-OO               C   8H  17O   2     G    300.00   3500.00 1600.00      1
 2.43863221e+01 4.79091863e-02-1.96116165e-05 3.85759153e-09-3.01446048e-13    2
-3.51809040e+04-9.31491997e+01-7.10506923e-01 1.10651259e-01-7.84323095e-05    3
 2.83662136e-08-4.13091825e-12-2.71499187e+04 3.97240936e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155885e+01 4.43694094e-02-1.35968858e-05 1.75327622e-09-6.83090880e-14    2
-3.76580614e+04-8.42148793e+01-5.96912081e+00 1.20872170e-01-9.61538217e-05    3
 4.13489289e-08-7.18982936e-12-3.02675122e+04 5.27954202e+01                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574275e-02-1.91478836e-05 3.78861311e-09-2.97862012e-13    2
-2.91331926e+04-1.00455337e+02-9.92411236e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
INDENE                  C   9H   8          G    300.00   3500.00 1450.00      1
 1.65348693e+01 2.81361431e-02-7.82674558e-06 2.33936401e-10 1.15234436e-13    2
 1.13278665e+04-6.66478053e+01-7.32592199e+00 9.39590155e-02-7.59193723e-05    3
 3.15408912e-08-5.28251639e-12 1.82474960e+04 5.73325203e+01                   4
INDENYL                 C   9H   7          G    300.00   3500.00 1600.00      1
 1.63412613e+01 3.01210631e-02-1.29067938e-05 2.63187626e-09-2.11554314e-13    2
 2.91054096e+04-6.81510017e+01-5.81714820e+00 8.55170869e-02-6.48405661e-05    3
 2.42709481e-08-3.59265929e-12 3.61961007e+04 4.91650485e+01                   4
KEA3B3                  C   3H   4O   4     G    300.00   3500.00 1500.00      1
 1.56495498e+01 1.47904715e-02-6.84032429e-06 1.49167145e-09-1.26830372e-13    2
-4.74213138e+04-4.92482738e+01 1.41905665e+00 5.27384532e-02-4.47883060e-05    3
 1.83574411e-08-2.93779198e-12-4.31521659e+04 2.51755980e+01                   4
KEA3G2                  C   3H   4O   4     G    300.00   3500.00 1540.00      1
 1.52972938e+01 1.47507483e-02-6.65907582e-06 1.42291765e-09-1.19027510e-13    2
-5.03228961e+04-4.71892678e+01 2.76516864e+00 4.73017226e-02-3.83645703e-05    3
 1.51482399e-08-2.34716424e-12-4.64630015e+04 1.86821429e+01                   4
KEHYBU1                 C   4H   8O   4     G    300.00   3500.00 1200.00      1
 1.50812003e+01 2.99746636e-02-1.37944087e-05 3.03171375e-09-2.60935208e-13    2
-6.34178095e+04-4.27051069e+01-4.53521777e+00 9.53627237e-02-9.55294839e-05    3
 4.84400888e-08-9.72101335e-12-5.87098692e+04 5.55092666e+01                   4
KEHYMB                  C   5H   8O   5     G    300.00   3500.00 1200.00      1
 1.28585854e+01 3.05267697e-02-1.05263784e-05 1.70287735e-09-1.06411281e-13    2
-6.04915273e+04-3.42459469e+01-2.28352158e+00 8.10004596e-02-7.36184908e-05    3
 3.67540509e-08-7.40873910e-12-5.68574216e+04 4.15666988e+01                   4
KHDECA                  C  10H  16O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415883e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853396e-05    3
 2.77298318e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   3500.00 1690.00      1
 6.18941987e+01 8.22994739e-02-3.10180668e-05 5.38913026e-09-3.62606874e-13    2
-9.79974660e+04-2.72277500e+02-3.09268744e+00 2.36114589e-01-1.67540358e-04    3
 5.92440776e-08-8.32931507e-12-7.60318984e+04 7.53471329e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076076e+01 1.68261952e-02-6.51181371e-06 1.21158891e-09-8.99428218e-14    2
 5.89425072e+04-3.55373248e+01 1.67614175e-01 5.94226632e-02-6.25597980e-05    3
 3.39881879e-08-7.27779348e-12 6.17104257e+04 2.46218079e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863876e+01 1.90072461e-02-7.30992558e-06 1.31482495e-09-9.21385789e-14    2
 3.55364843e+04-4.09021933e+01-1.05889383e+00 6.36321466e-02-6.08598062e-05    3
 2.98747613e-08-5.80412585e-12 3.90228046e+04 2.94875281e+01                   4
MACRIL                  C   4H   6O   2     G    300.00   3500.00 1110.00      1
 9.14034166e+00 2.10870489e-02-7.42259222e-06 1.25044332e-09-8.33064060e-14    2
-4.12827789e+04-1.50267978e+01-1.13135763e+00 5.81021815e-02-5.74430417e-05    3
 3.12927553e-08-6.84959289e-12-3.90024617e+04 3.56001684e+01                   4
MB                      C   5H  10O   2     G    300.00   3500.00 1800.00      1
 1.24284224e+01 3.57133446e-02-1.61592883e-05 3.52094113e-09-3.02693515e-13    2
-6.07702348e+04-3.65220690e+01 2.77831320e+00 5.71580318e-02-3.40298609e-05    3
 1.01396717e-08-1.22196165e-12-5.72961955e+04 1.57063351e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1540.00      1
 1.14154101e+01 2.70830264e-02-1.13419491e-05 2.30157826e-09-1.86056675e-13    2
 6.23040748e+03-4.10347479e+01-6.52219774e+00 7.36742157e-02-5.67229776e-05    3
 2.19470452e-08-3.37525585e-12 1.17551907e+04 5.32489849e+01                   4
MCROT                   C   5H   8O   2     G    300.00   3500.00 1270.00      1
 1.13738847e+01 2.61318034e-02-8.74855171e-06 1.35831508e-09-8.00175020e-14    2
-4.63062146e+04-2.54801461e+01 2.72064727e-01 6.10981657e-02-5.00474047e-05    3
 2.30375030e-08-4.34757418e-12-4.34863523e+04 3.07332406e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194568e+01 4.36180644e-02-1.87773363e-05 3.92059023e-09-3.26702984e-13    2
-2.91866300e+04-7.40611877e+01-1.01006358e+01 1.03218270e-01-6.84441744e-05    3
 2.23157154e-08-2.88158149e-12-1.95313967e+04 7.10947481e+01                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317081e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
MCYC6-OQOOH             C   7H  12O   3     G    300.00   3500.00 1800.00      1
 2.89245833e+01 2.89702632e-02-1.00807411e-05 1.60861341e-09-9.81376976e-14    2
-5.92858085e+04-1.29605491e+02-5.14358533e+00 1.04677305e-01-7.31699422e-05    3
 2.49749842e-08-3.34346697e-12-4.70212678e+04 5.47785441e+01                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522001e-06 1.12153176e-09-5.23348938e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317081e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522001e-06 1.12153176e-09-5.23348938e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MD                      C  11H  22O   2     G    300.00   3500.00 1800.00      1
 3.32942906e+01 6.02278032e-02-2.43433721e-05 4.77523421e-09-3.75629873e-13    2
-8.61538195e+04-1.40508531e+02 1.40263274e+00 1.31098154e-01-8.34019977e-05    3
 2.66487992e-08-3.41362502e-12-7.46728226e+04 3.20957740e+01                   4
MDKETO                  C  11H  20O   5     G    300.00   3500.00 1420.00      1
 2.98411867e+01 7.16595718e-02-3.12595573e-05 6.71204593e-09-5.73522120e-13    2
-1.08207342e+05-1.07784039e+02 3.72296254e+00 1.45232034e-01-1.08976947e-04    3
 4.31990835e-08-6.99729634e-12-1.00789766e+05 2.73798301e+01                   4
MEFU2                   C   5H   6O   1     G    300.00   3500.00 1260.00      1
 5.16398169e+00 3.29529080e-02-1.68209195e-05 4.03716052e-09-3.55511369e-13    2
-1.31841670e+04-2.67616710e+00-3.74149804e+00 6.12242723e-02-5.04773055e-05    3
 2.18447722e-08-3.88876765e-12-1.09399861e+04 4.23457855e+01                   4
MEK                     C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.00996674e+01 2.22850926e-02-8.24112797e-06 1.42760366e-09-9.77654881e-14    2
-3.40270944e+04-2.55002808e+01 1.67138626e+00 4.10146063e-02-2.38490560e-05    3
 7.20831776e-09-9.00642446e-13-3.09929132e+04 2.01153350e+01                   4
MEOLE                   C  19H  36O   2     G    300.00   3500.00 1800.00      1
 5.99431010e+01 8.58698597e-02-2.97675970e-05 4.64267973e-09-2.70021412e-13    2
-1.05323856e+05-2.71321378e+02-2.40342610e-02 2.19130160e-01-1.40817847e-04    3
 4.57724021e-08-5.98248285e-12-8.37356873e+04 5.32332675e+01                   4
MLIN1                   C  19H  32O   2     G    300.00   3500.00 1790.00      1
 6.02396272e+01 7.58944997e-02-2.57645248e-05 3.83449043e-09-2.03418185e-13    2
-7.74468689e+04-2.75096818e+02-2.53501097e+00 2.16173021e-01-1.43316358e-04    3
 4.76154339e-08-6.31807509e-12-5.49735485e+04 6.43028989e+01                   4
MLINO                   C  19H  34O   2     G    300.00   3500.00 1800.00      1
 6.05955674e+01 8.00185064e-02-2.72219227e-05 4.09057977e-09-2.22036540e-13    2
-9.16175365e+04-2.76065905e+02-1.22142744e+00 2.17389606e-01-1.41697839e-04    3
 4.64890673e-08-6.11071537e-12-6.93634183e+04 5.85005668e+01                   4
MPA                     C  17H  34O   2     G    300.00   3500.00 1570.00      1
 4.76347765e+01 8.91363271e-02-3.14080949e-05 4.73916072e-09-2.33379401e-13    2
-1.08404908e+05-2.13800451e+02-6.71212905e+00 2.27599781e-01-1.63698019e-04    3
 6.09132260e-08-9.17829426e-12-9.13399797e+04 7.29065166e+01                   4
MSTEA                   C  19H  38O   2     G    300.00   3500.00 1590.00      1
 5.57521885e+01 9.44092844e-02-3.21197984e-05 4.65296638e-09-2.12922185e-13    2
-1.17225837e+05-2.54579461e+02-7.52353560e+00 2.53593496e-01-1.82293583e-04    3
 6.76189138e-08-1.01132284e-11-9.71041567e+04 8.00324369e+01                   4
MSTEAKETO               C  19H  36O   5     G    300.00   3500.00 1630.00      1
 6.13348222e+01 9.80436966e-02-3.77033724e-05 6.80817282e-09-4.83388457e-13    2
-1.42870185e+05-2.70834349e+02-4.17722454e-01 2.49583683e-01-1.77157348e-04    3
 6.38445637e-08-9.23130116e-12-1.22738855e+05 5.72570421e+01                   4
MTBE                    C   5H  12O   1     G    300.00   3500.00 1320.00      1
 9.85250854e+00 4.01896195e-02-1.66704212e-05 3.10158953e-09-2.11537799e-13    2
-4.09274217e+04-2.61941109e+01-1.85856423e+00 7.56777188e-02-5.69978068e-05    3
 2.34689560e-08-4.06899357e-12-3.78356985e+04 3.35564110e+01                   4
MTBE-O                  C   5H  10O   2     G    300.00   3500.00 1520.00      1
 1.51388759e+01 2.99979380e-02-1.22799224e-05 2.46100800e-09-1.97690794e-13    2
-5.39879921e+04-5.57113238e+01-5.03717524e+00 8.30928094e-02-6.46761770e-05    3
 2.54418214e-08-3.97742985e-12-4.78544725e+04 5.00743811e+01                   4
MTBE-OO                 C   5H  11O   3     G    300.00   3500.00 1650.00      1
 1.64806404e+01 3.48147986e-02-1.47688716e-05 3.00165535e-09-2.41352124e-13    2
-3.59678540e+04-5.02874924e+01 2.84930352e+00 6.78604638e-02-4.48103854e-05    3
 1.51396407e-08-2.08044082e-12-3.14695128e+04 2.23020650e+01                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   3500.00 1360.00      1
 1.70053287e+01 4.31260455e-02-1.99573148e-05 4.44658587e-09-3.89314847e-13    2
-4.64302952e+04-4.61328184e+01 4.65469152e+00 7.94514489e-02-6.00220979e-05    3
 2.40861854e-08-3.99953536e-12-4.30709219e+04 1.72494984e+01                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   3500.00 1750.00      1
 2.60727575e+01 2.16561735e-02-7.50837024e-06 1.18094191e-09-6.95946679e-14    2
-6.60762157e+04-1.03020582e+02 2.39248713e+00 7.57825058e-02-5.39023694e-05    3
 1.88548464e-08-2.59443816e-12-5.77881211e+04 2.44748876e+01                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   3500.00 1320.00      1
 1.54436171e+01 3.66620452e-02-1.53964703e-05 3.18866664e-09-2.64826209e-13    2
-2.86187067e+04-4.25445321e+01 1.39866729e+00 7.92224991e-02-6.37606224e-05    3
 2.76150061e-08-4.89102686e-12-2.49108399e+04 2.91135557e+01                   4
N                       N   1               G    300.00   3500.00 1800.00      1
 2.43583682e+00 1.27743369e-04-8.58132365e-08 2.13268140e-11-1.23433516e-15    2
 5.61236145e+04 4.53259076e+00 2.50515554e+00-2.62982346e-05 4.25547663e-08    3
-2.62168907e-11 5.36895716e-15 5.60986597e+04 4.15742338e+00                   4
N1C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.19078661e+01 2.67959929e-02-1.07944841e-05 2.10106148e-09-1.63536607e-13    2
-3.95221179e+04-3.57389868e+01 7.73360084e-02 5.30860597e-02-3.27028730e-05    3
 1.02152796e-08-1.29051135e-12-3.52631271e+04 2.82903098e+01                   4
N2                      N   2               G    300.00   3500.00 1050.00      1
 2.71287897e+00 1.90359754e-03-8.54297556e-07 1.84170938e-10-1.54715988e-14    2
-8.40225273e+02 7.15926558e+00 3.85321336e+00-2.44053349e-03 5.35160392e-06    3
-3.75608397e-09 9.22684330e-13-1.07969550e+03 1.60217419e+00                   4
N2C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.39850075e+01 2.35768220e-02-8.73106106e-06 1.51546163e-09-1.02847459e-13    2
-4.24053999e+04-4.83702850e+01 1.11912948e-01 5.44059211e-02-3.44219770e-05    3
 1.10306157e-08-1.42439663e-12-3.74110858e+04 2.67137970e+01                   4
N2H2                    H   2N   2          G    300.00   3500.00  930.00      1
 1.94872574e+00 9.02206572e-03-4.48167913e-06 1.07159624e-09-9.96387287e-14    2
 2.46850174e+04 1.27074554e+01 2.44745784e+00 6.87698140e-03-1.02186571e-06    3
-1.40855675e-09 5.67069064e-13 2.45922533e+04 1.03375547e+01                   4
N2H3                    H   3N   2          G    300.00   3500.00 1610.00      1
 5.06961797e+00 6.18061831e-03-1.87909018e-06 2.33273638e-10-8.03110073e-15    2
 1.63477734e+04-4.00218491e+00 1.71415249e+00 1.45171785e-02-9.64607174e-06    3
 3.44941507e-09-5.07431944e-13 1.74282333e+04 1.37839838e+01                   4
N2H4                    H   4N   2          G    300.00   3500.00 1160.00      1
 4.91914378e+00 9.71187969e-03-3.62925367e-06 6.36530934e-10-4.28508947e-14    2
 9.36304606e+03-2.64395648e+00 3.60425651e-01 2.54315974e-02-2.39564748e-05    3
 1.23188419e-08-2.56059034e-12 1.04206687e+04 2.00258283e+01                   4
N2O                     O   1N   2          G    300.00   3500.00 1650.00      1
 5.52129143e+00 1.46645965e-03-3.04694075e-07-1.87106858e-11 8.50389041e-15    2
 7.81312268e+03-6.17451657e+00 2.68521969e+00 8.34178508e-03-6.55498992e-06    3
 2.50666137e-09-3.74128239e-13 8.74902635e+03 8.92812480e+00                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   3500.00 1800.00      1
 4.08087723e+01 4.96339543e-02-1.81420129e-05 3.12006732e-09-2.11175642e-13    2
-5.65432959e+04-1.73811020e+02 2.62701325e+00 1.34482308e-01-8.88489740e-05    3
 2.93078307e-08-3.84836500e-12-4.27978627e+04 3.28366249e+01                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   3500.00 1650.00      1
 2.99089271e+01 5.87016386e-02-2.37959516e-05 4.63914804e-09-3.59659107e-13    2
-7.07246459e+04-1.14602343e+02 2.87865509e+00 1.24229571e-01-8.33667990e-05    3
 2.87081773e-08-4.00648172e-12-6.18046561e+04 2.93391873e+01                   4
NC10-QOOH               C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.67714538e+01 4.56787199e-02-1.56929249e-05 2.49979255e-09-1.53467299e-13    2
-3.72897414e+04-1.54708984e+02 8.46533635e-01 1.25511876e-01-8.22205548e-05    3
 2.71396555e-08-3.57567048e-12-2.43567701e+04 3.97241784e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971791e+01 4.89478938e-02-1.82737062e-05 3.23575201e-09-2.26811843e-13    2
-3.12534582e+04-1.16784058e+02-2.31417710e+00 1.16973130e-01-7.49614029e-05    3
 2.42311952e-08-3.14284562e-12-2.02333700e+04 4.88909878e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212692e+01 5.52219738e-02-2.21266526e-05 4.33498891e-09-3.42316503e-13    2
-2.10175171e+04-1.03192977e+02-1.81057271e+00 1.17737178e-01-7.42226562e-05    3
 2.36298050e-08-3.02215208e-12-1.08900540e+04 4.90624204e+01                   4
NC10H21-OO              C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.23779830e+01 5.24885367e-02-1.93370131e-05 3.35369674e-09-2.28448799e-13    2
-4.06447276e+04-1.32098961e+02 1.67478189e+00 1.20717872e-01-7.61947929e-05    3
 2.44121337e-08-3.15323171e-12-2.95915752e+04 3.40731686e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878918e+01 5.29920990e-02-1.98404553e-05 3.55616370e-09-2.54281184e-13    2
-4.56232379e+04-1.22752047e+02-2.17870143e+00 1.22917862e-01-7.81119243e-05    3
 2.51381893e-08-3.25178473e-12-3.42952643e+04 4.75517200e+01                   4
NC10MOOH                C  10H  20O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889668e+01 5.84439691e-02-2.09491580e-05 3.49897609e-09-2.27324946e-13    2
-6.45487872e+04-2.03262107e+02 2.75932352e+00 1.56509843e-01-1.02670720e-04    3
 3.37662211e-08-4.43110898e-12-4.86621157e+04 3.55767286e+01                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762540e+01 8.51935060e-02-4.32222039e-05 1.03184896e-08-9.52873634e-13    2
-7.66784457e+04-1.07151303e+02 4.95723376e+00 1.38569107e-01-8.77018710e-05    3
 2.67924404e-08-3.24092235e-12-6.80315984e+04 2.28446447e+01                   4
NC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763735e+01 5.51011626e-02-1.90602563e-05 3.05791504e-09-1.89217484e-13    2
-4.53973988e+04-1.84606456e+02 5.27389362e-01 1.49210016e-01-9.74843011e-05    3
 3.21038575e-08-4.22337617e-12-3.01517645e+04 4.45950809e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295229e-05 5.21804509e-09-4.10998518e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710595e-12-1.66984825e+04 5.11161660e+01                   4
NC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754174e+01 6.23046009e-02-2.29785783e-05 3.99220438e-09-2.72630412e-13    2
-4.86703034e+04-1.60846136e+02 1.39669302e+00 1.44257322e-01-9.12725124e-05    3
 2.92862540e-08-3.78569287e-12-3.53939626e+04 3.87492139e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414095e+01 6.11045883e-02-2.24641073e-05 3.93182440e-09-2.73349362e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1800.00      1
 5.83925916e+01 7.87490301e-02-2.86987240e-05 4.90944000e-09-3.29403315e-13    2
-8.05061539e+04-2.59209019e+02 2.14519035e+00 2.03743255e-01-1.32860578e-04    3
 4.34879045e-08-5.68752339e-12-6.02570894e+04 4.52136503e+01                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1690.00      1
 4.88441297e+01 8.47833151e-02-3.17577492e-05 5.56702742e-09-3.82331487e-13    2
-9.50808904e+04-2.07202631e+02 1.75040694e+00 1.96247748e-01-1.30690678e-04    3
 4.45938236e-08-6.15552619e-12-7.91632121e+04 4.47087787e+01                   4
NC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.49634696e+01 7.74662171e-02-2.71265902e-05 4.36953904e-09-2.68719606e-13    2
-8.49949222e+04-2.46825964e+02 8.02842616e-02 1.99428851e-01-1.28762119e-04    3
 4.20123273e-08-5.49688464e-12-6.52369755e+04 5.02132837e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278372e+01 8.00212238e-02-3.03236333e-05 5.55903616e-09-4.09822553e-13    2
-4.61545210e+04-2.04019481e+02-3.22413374e+00 1.90803381e-01-1.22642098e-04    3
 3.97510601e-08-5.15871477e-12-2.82078115e+04 6.57897858e+01                   4
NC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.00344484e+01 8.20070153e-02-3.03042993e-05 5.28016700e-09-3.62022840e-13    2
-6.47045872e+04-2.18137205e+02 8.65096715e-01 1.91272241e-01-1.21358654e-04    3
 3.90040022e-08-5.04588884e-12-4.70036206e+04 4.79775838e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210237e+01 7.73881688e-02-2.77557896e-05 4.69678103e-09-3.12959243e-13    2
-7.08514664e+04-2.24842855e+02-3.64057977e+00 1.96191732e-01-1.26758759e-04    3
 4.13645475e-08-5.40570458e-12-5.16052891e+04 6.45024955e+01                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1260.00      1
 1.11683562e+01 2.95822139e-02-1.42526305e-05 3.27126849e-09-2.92476812e-13    2
-2.00281219e+04-2.06289848e+01 2.57588692e+00 5.68598942e-02-4.67260594e-05    3
 2.04529769e-08-3.70154594e-12-1.78628196e+04 2.28105329e+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1800.00      1
 1.29748618e+01 1.76433870e-02-7.16935406e-06 1.42696153e-09-1.14477043e-13    2
-5.86411825e+03-3.67690498e+01 1.55643299e+00 4.30176732e-02-2.83145926e-05    3
 9.25853134e-09-1.20219507e-12-1.75348388e+03 2.50298688e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1650.00      1
 8.44692954e+00 1.52881013e-02-4.72394213e-06 3.72053769e-10 2.77825399e-14    2
 7.24499466e+03-1.97652064e+01 5.40130268e-01 3.44560996e-02-2.21493951e-05    3
 7.41264082e-09-1.03897307e-12 9.85423842e+03 2.23400592e+01                   4
NC3H7O                  C   3H   7O   1     G    300.00   3500.00 1800.00      1
 9.66226461e+00 1.80582994e-02-6.80752580e-06 1.22634214e-09-8.79552073e-14    2
-9.72942766e+03-2.55365895e+01-5.52121379e-01 4.07569349e-02-2.57230554e-05    3
 8.23209384e-09-1.06097628e-12-6.05224870e+03 2.97457983e+01                   4
NC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1800.00      1
 1.03578665e+01 1.87834500e-02-6.54155125e-06 1.06792692e-09-6.79101580e-14    2
-3.60054458e+04-2.89224528e+01 2.34636347e-01 4.12795171e-02-2.52882738e-05    3
 8.01115750e-09-1.03224774e-12-3.23610829e+04 2.58665808e+01                   4
NC3H7OO                 C   3H   7O   2     G    300.00   3500.00 1650.00      1
 9.25591855e+00 2.27563801e-02-9.54934453e-06 1.92559464e-09-1.53946670e-13    2
-9.34005086e+03-1.86388081e+01 1.92964396e+00 4.05170458e-02-2.56954042e-05    3
 8.44925513e-09-1.14238008e-12-6.92238025e+03 2.03750491e+01                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   3500.00 1230.00      1
 1.51474113e+01 3.37812811e-02-1.58996825e-05 3.57608795e-09-3.14486517e-13    2
-2.85698876e+04-4.24732203e+01 1.10123476e+00 7.94599040e-02-7.16053202e-05    3
 3.37688455e-08-6.45122586e-12-2.51145282e+04 2.81992197e+01                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1330.00      1
 1.18153445e+01 3.20093755e-02-1.53334981e-05 3.50316407e-09-3.12136547e-13    2
-4.27660549e+04-2.73083214e+01 2.51946600e+00 5.99669047e-02-4.68645461e-05    3
 1.93082006e-08-3.28300808e-12-4.02933512e+04 2.01899074e+01                   4
NC4-QOOH                C   4H   9O   2     G    300.00   3500.00 1760.00      1
 1.83774568e+01 1.83354725e-02-6.23923380e-06 9.66797421e-10-5.61281943e-14    2
-1.29135491e+04-6.55986639e+01 1.19976578e+00 5.73756794e-02-3.95121374e-05    3
 1.35701700e-08-1.84637998e-12-6.86700189e+03 2.69845517e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14852000e-06-5.94424182e-11 5.32964635e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
NC4H8                   C   4H   8          G    300.00   3500.00 1170.00      1
 2.98709814e+00 3.25282541e-02-1.46250479e-05 2.94136385e-09-2.14960813e-13    2
-2.50111901e+03 1.03971909e+01-1.05707773e+00 4.63544964e-02-3.23509995e-05    3
 1.30416212e-08-2.37313546e-12-1.55478186e+03 3.05429525e+01                   4
NC4H9-OO                C   4H   9O   2     G    300.00   3500.00 1320.00      1
 8.96630114e+00 3.41074657e-02-1.57641000e-05 3.50715782e-09-3.06662916e-13    2
-1.40847395e+04-1.58347447e+01 9.44281655e-01 5.84166156e-02-4.33881341e-05    3
 1.74586902e-08-2.94899859e-12-1.19669263e+04 2.50940293e+01                   4
NC4H9P                  C   4H   9          G    300.00   3500.00  950.00      1
 3.94763005e+00 3.16286394e-02-1.12984867e-05 1.11637452e-09 5.54031592e-14    2
 6.05554723e+03 7.76350069e+00-2.76188363e-01 4.94131380e-02-3.93792739e-05    3
 2.08221901e-08-5.13033778e-12 6.85807273e+03 2.79243294e+01                   4
NC4H9S                  C   4H   9          G    300.00   3500.00  850.00      1
 3.40122925e+00 3.20901864e-02-1.12255471e-05 9.71712129e-10 8.30726251e-14    2
 4.66283102e+03 1.05291640e+01 2.36336476e-01 4.69837994e-02-3.75083937e-05    3
 2.15857094e-08-5.97986776e-12 5.20086279e+03 2.52835872e+01                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   3500.00 1270.00      1
 1.54638476e+01 4.30531975e-02-2.04284728e-05 4.63174721e-09-4.10271992e-13    2
-3.17413365e+04-4.31406917e+01 1.43265566e+00 8.72459280e-02-7.26246113e-05    3
 3.20312950e-08-5.80388375e-12-2.81774138e+04 2.79053907e+01                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   3500.00 1410.00      1
 1.42172630e+01 3.77707683e-02-1.76257936e-05 3.93443034e-09-3.43954252e-13    2
-4.65061050e+04-3.85369191e+01 2.52749929e+00 7.09332187e-02-5.29049961e-05    3
 2.06149043e-08-3.30148510e-12-4.32095916e+04 2.18759162e+01                   4
NC5-QOOH                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.36538194e+01 3.77860020e-02-1.75151081e-05 3.90394425e-09-3.41708560e-13    2
-1.43879859e+04-3.94678819e+01-5.74283055e-01 8.15647789e-02-6.80290814e-05    3
 2.98085460e-08-5.32336273e-12-1.06886793e+04 3.29074336e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929736e+01 2.82582223e-02-1.13863841e-05 2.22526491e-09-1.74280993e-13    2
-1.02483443e+04-3.39253533e+01-6.89551964e-01 5.46638348e-02-3.33910611e-05    3
 1.03751453e-08-1.30620882e-12-5.97063504e+03 3.03853541e+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.40073101e+01 3.04405284e-02-1.35854526e-05 2.90305354e-09-2.44985844e-13    2
-2.55455866e+04-5.25239383e+01-3.79263098e+00 6.99959530e-02-4.65483064e-05    3
 1.51115179e-08-1.94060590e-12-1.91376078e+04 4.38130562e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93193785e+00 3.75440987e-02-1.65478566e-05 3.53633643e-09-2.99976701e-13    2
-1.73087074e+03-8.88710670e+00-3.57520449e+00 6.08933039e-02-3.60055276e-05    3
 1.07428812e-08-1.30088570e-12 2.05170050e+03 4.79797395e+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   3500.00 1630.00      1
 1.66988185e+01 3.44172712e-02-1.43139761e-05 2.85300849e-09-2.25350876e-13    2
-3.73755763e+04-5.75775303e+01 6.24289371e-02 7.52427671e-02-5.18834508e-05    3
 1.82188468e-08-2.58207455e-12-3.19521133e+04 3.08116402e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559082e+01 1.49866375e-02-1.56738312e-06-4.84518435e-10 9.00436509e-14    2
-2.80668702e+04-9.05497671e+01-1.97000865e+00 6.65997861e-02-4.45783403e-05    3
 1.54454657e-08-2.12245414e-12-1.97055401e+04 3.51537401e+01                   4
NC5H12OO                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.06544848e+01 4.16170555e-02-1.93382868e-05 4.32113942e-09-3.79088223e-13    2
-1.98652039e+04-2.50234586e+01 3.19664880e-01 7.34165014e-02-5.60299551e-05    3
 2.31373796e-08-3.99759595e-12-1.71781508e+04 2.75475609e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951654e+01 5.24635942e-03 6.43208138e-06-3.19131389e-09 4.01093698e-13    2
-1.79767847e+04-1.24497292e+02-1.85358315e+00 7.25469181e-02-5.02818725e-05    3
 1.80498673e-08-2.58221827e-12-7.31503024e+03 3.72569567e+01                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   3500.00 1690.00      1
 2.24694069e+01 4.29307086e-02-1.68910162e-05 3.18431082e-09-2.38592446e-13    2
-4.58962940e+04-7.93472401e+01 2.87430503e+00 8.93096479e-02-5.80557552e-05    3
 1.94228666e-08-2.64074567e-12-3.92731495e+04 2.54699082e+01                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   3500.00 1670.00      1
 2.27584121e+01 4.25741258e-02-1.77950010e-05 3.55398722e-09-2.80791799e-13    2
-5.95329656e+04-8.19251639e+01 2.24997334e+00 9.16961348e-02-6.19165660e-05    3
 2.11673864e-08-2.91752820e-12-5.26831470e+04 2.75334100e+01                   4
NC7-QOOH                C   7H  15O   2     G    300.00   3500.00 1800.00      1
 3.67777501e+01 2.43465392e-02-1.65378817e-05 5.22869888e-09-5.85107382e-13    2
-2.84549794e+04-1.65059640e+02-2.87358792e+00 1.12460624e-01-8.99662853e-05    3
 3.24244039e-08-4.36228864e-12-1.41804977e+04 4.95416730e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360661e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC7H13OOH               C   7H  14O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668105e+01 3.59607890e-02-1.37346402e-05 2.52229050e-09-1.85248240e-13    2
-1.87497345e+04-6.92309265e+01-1.22797309e+00 7.92825302e-02-4.98360912e-05    3
 1.58931983e-08-2.04231877e-12-1.17316124e+04 3.62789089e+01                   4
NC7H14O                 C   7H  14O   1     G    300.00   3500.00 1490.00      1
 1.37609323e+01 4.99379374e-02-2.21152348e-05 4.72010363e-09-3.98160014e-13    2
-3.97917916e+04-4.67908592e+01-7.39181743e+00 1.06723843e-01-7.92822536e-05    3
 3.02981881e-08-4.68978493e-12-3.34882722e+04 6.36941424e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938298e+01 4.32851195e-02-1.83429598e-05 3.81524632e-09-3.18291961e-13    2
-8.33589206e+03-5.34387877e+01-1.03213606e+00 8.08983770e-02-4.96873411e-05    3
 1.54242764e-08-1.93065725e-12-2.24254435e+03 3.81680705e+01                   4
NC7H15-OO               C   7H  15O   2     G    300.00   3500.00 1780.00      1
 2.68006146e+01 3.35780866e-02-1.17982179e-05 1.89992229e-09-1.16218734e-13    2
-2.33388920e+04-1.06550436e+02 1.92333992e+00 8.94820746e-02-5.89083201e-05    3
 1.95441553e-08-2.59434135e-12-1.44825822e+04 2.78126029e+01                   4
NC7H15OOH               C   7H  16O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696120e+01 1.73458864e-02-4.57663884e-07-1.06280964e-09 1.59098857e-13    2
-3.76541592e+04-1.40920497e+02-2.76912812e+00 9.25430866e-02-6.31219974e-05    3
 2.21462028e-08-3.06437509e-12-2.54722127e+04 4.22218230e+01                   4
NCO                     C   1O   1N   1     G    300.00   3500.00 1700.00      1
 5.80612871e+00 1.29457396e-03-2.96387145e-07-4.45669057e-12 6.00806513e-15    2
 1.70053704e+04-6.33800183e+00 2.87969597e+00 8.18029805e-03-6.37202605e-06    3
 2.37814680e-09-3.44374801e-13 1.80003575e+04 9.33319238e+00                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   3500.00 1800.00      1
 2.53088279e+01 2.46008468e-02-8.38584870e-06 1.28446216e-09-7.25492020e-14    2
-3.52662111e+04-9.88693150e+01 2.93992987e+00 7.43095092e-02-4.98097340e-05    3
 1.66266419e-08-2.20340750e-12-2.72134078e+04 2.21958278e+01                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   3500.00 1690.00      1
 2.24459936e+01 2.37621277e-02-8.83881473e-06 1.53830075e-09-1.04514815e-13    2
-5.03880249e+04-8.77405631e+01 1.27283562e+00 7.38761111e-02-5.33186817e-05    3
 1.90845993e-08-2.70012112e-12-4.32314975e+04 2.55178450e+01                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   3500.00 1630.00      1
 1.86197530e+01 2.85111424e-02-1.13969334e-05 2.18137254e-09-1.65768942e-13    2
-1.50391446e+04-6.74883738e+01 1.48070310e+00 7.05701605e-02-5.01015514e-05    3
 1.80114821e-08-2.59369986e-12-9.45181437e+03 2.35714319e+01                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   3500.00 1470.00      1
 1.29296103e+01 3.16150611e-02-1.35584975e-05 2.81753187e-09-2.32686285e-13    2
-2.37933924e+04-4.88968548e+01-6.91462638e+00 8.56129839e-02-6.86584188e-05    3
 2.78061583e-08-4.48245268e-12-1.79591868e+04 5.44853542e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276289e+01 2.66845577e-02-1.02158264e-05 1.86929104e-09-1.35803312e-13    2
-2.94216421e+03-5.15145769e+01-1.29689709e+00 6.41085720e-02-4.38302105e-05    3
 1.52882069e-08-2.14462305e-12 2.27642747e+03 3.18773552e+01                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   3500.00 1660.00      1
 1.69989732e+01 3.01601499e-02-1.19254896e-05 2.25822367e-09-1.69878947e-13    2
-2.10464569e+04-6.14617731e+01 1.07910948e+00 6.85212672e-02-4.65891499e-05    3
 1.61793724e-08-2.26643749e-12-1.57610621e+04 2.34108339e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220811e+01 2.73824077e-02-1.01392581e-05 1.77707009e-09-1.22756971e-13    2
-2.85197010e+04-6.62488521e+01-2.62463460e+00 7.07864446e-02-4.84369376e-05    3
 1.67957680e-08-2.33138901e-12-2.22478177e+04 3.25342362e+01                   4
NH                      H   1N   1          G    300.00   3500.00 1550.00      1
 2.53691464e+00 1.74532708e-03-6.66818142e-07 1.34160653e-10-1.04190033e-14    2
 4.21821879e+04 7.12732805e+00 3.75007687e+00-1.38541418e-03 2.36293147e-06    3
-1.16895746e-09 1.99761337e-13 4.18061076e+04 7.42847188e-01                   4
NH2                     H   2N   1          G    300.00   3500.00 1120.00      1
 2.67687765e+00 3.48484078e-03-1.28570820e-06 2.72091630e-10-2.36034281e-14    2
 2.20303372e+04 7.34730162e+00 4.18313061e+00-1.89463407e-03 5.91894562e-06    3
-4.01639279e-09 9.33647558e-13 2.16929365e+04-9.01998745e-02                   4
NH3                     H   3N   1          G    300.00   3500.00 1210.00      1
 2.21117984e+00 6.52182453e-03-2.30931532e-06 3.98907128e-10-2.80385645e-14    2
-6.39009604e+03 8.86905603e+00 3.21689186e+00 3.19715670e-03 1.81217371e-06    3
-1.87188573e-09 4.41133513e-13-6.63347835e+03 3.82536772e+00                   4
NNH                     H   1N   2          G    300.00   3500.00  720.00      1
 2.67540125e+00 5.35668680e-03-2.94990450e-06 7.78541240e-10-7.91413867e-14    2
 2.84746064e+04 1.03028707e+01 3.96823590e+00-1.82572793e-03 1.20134595e-05    3
-1.30764254e-08 4.73161093e-12 2.82884383e+04 4.49039228e+00                   4
NO                      O   1N   1          G    300.00   3500.00  970.00      1
 2.69775018e+00 2.39887133e-03-1.31644700e-06 3.38235813e-10-3.29394890e-14    2
 9.99854348e+03 9.40230813e+00 3.91290193e+00-2.61206371e-03 6.43242163e-06    3
-4.98744709e-09 1.33965920e-12 9.76280404e+03 3.57691592e+00                   4
NO2                     O   2N   1          G    300.00   3500.00 1800.00      1
 5.25673685e+00 1.64343307e-03-6.24197948e-07 1.07065150e-10-6.88584753e-15    2
 1.95363563e+03-2.35827568e+00 2.61409592e+00 7.51596848e-03-5.51797745e-06    3
 1.91957608e-09-2.58623476e-13 2.90498637e+03 1.19442483e+01                   4
NO3                     O   3N   1          G    300.00   3500.00 1330.00      1
 7.66391925e+00 2.28165967e-03-8.16241554e-07 1.11367864e-10-3.38429715e-15    2
 5.62975022e+03-1.51899442e+01 4.06541943e-01 2.41083583e-02-2.54328190e-05    3
 1.24505044e-08-2.32277087e-12 7.56021258e+03 2.18923574e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963371e+01 3.80090295e-02-1.52789389e-05 2.95630099e-09-2.27699217e-13    2
-8.96605283e+03-7.62711275e+01-5.58650157e+00 9.92161261e-02-7.26605920e-05    3
 2.68653231e-08-3.96348393e-12-1.13154446e+03 5.33514397e+01                   4
O                       O   1               G    300.00   3500.00  950.00      1
 2.57318360e+00-8.95609984e-05 4.05096303e-08-8.39812674e-12 9.43621991e-16    2
 2.92191409e+04 4.74952023e+00 2.95200330e+00-1.68459131e-03 2.55897854e-06    3
-1.77574473e-09 4.66034833e-13 2.91471652e+04 2.94136507e+00                   4
O2                      O   2               G    300.00   3500.00  760.00      1
 2.81750648e+00 2.49838007e-03-1.52493521e-06 4.50547608e-10-4.87702792e-14    2
-9.31713392e+02 7.94729337e+00 3.46035080e+00-8.85011121e-04 5.15281056e-06    3
-5.40712413e-09 1.87809542e-12-1.02942573e+03 5.02236126e+00                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109941e+01 4.74108396e-02-1.82963852e-05 3.42084161e-09-2.57817125e-13    2
-2.68355230e+04-1.31410203e+02-1.02710769e+01 1.32926553e-01-8.95594797e-05    3
 2.98145803e-08-3.92361417e-12-1.29819774e+04 7.68627930e+01                   4
OH                      H   1O   1          G    300.00   3500.00  880.00      1
 3.62538436e+00-5.02165281e-04 8.36958463e-07-2.95714531e-10 3.30350486e-14    2
 3.41380110e+03 1.55419440e+00 3.37995109e+00 6.13440526e-04-1.06464235e-06    3
 1.14489214e-09-3.76228211e-13 3.45699735e+03 2.70689352e+00                   4
PC3H4                   C   3H   4          G    300.00   3500.00  920.00      1
 3.04156590e+00 1.80732925e-02-9.19849468e-06 2.29161583e-09-2.25689445e-13    2
 2.06214251e+04 7.37493873e+00 1.35943188e+00 2.53869187e-02-2.11228852e-05    3
 1.09324785e-08-2.57374996e-12 2.09309378e+04 1.53500040e+01                   4
QBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1270.00      1
 9.44680463e+00 1.40890825e-02-6.70668585e-06 1.51288685e-09-1.32818576e-13    2
 1.91332917e+04-2.81812927e+01-5.88861871e+00 6.23896285e-02-6.37545748e-05    3
 3.14592852e-08-6.02777889e-12 2.30284892e+04 4.94686856e+01                   4
QDECOOH                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
QMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557066e+01 1.60203243e-02-2.33018024e-06-2.09432791e-10 5.96256606e-14    2
-5.87318865e+04-9.28197844e+01-3.02577545e+00 9.80395304e-02-9.34626315e-05    3
 4.47942468e-08-8.27438909e-12-5.12578864e+04 4.90347050e+01                   4
QMDOOH                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.77681786e+01 6.05584838e-02-2.66377343e-05 5.63139231e-09-4.71383628e-13    2
-7.68263296e+04-1.55143375e+02 4.12866858e+00 1.35312950e-01-8.89331232e-05    3
 2.87037586e-08-3.67587894e-12-6.47161060e+04 2.69206708e+01                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 6.66288425e+01 8.44466273e-02-2.89700155e-05 4.40900507e-09-2.44932292e-13    2
-1.50877986e+05-3.00442019e+02-9.98790182e-01 2.34730256e-01-1.54206372e-04    3
 5.07928409e-08-6.68713172e-12-1.26532038e+05 6.55728373e+01                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1610.00      1
 5.66825541e+01 9.03049166e-02-3.59434818e-05 6.72610917e-09-4.95506768e-13    2
-6.74923687e+04-2.44601780e+02-2.71828911e+00 2.37884651e-01-1.73440129e-04    3
 6.36605386e-08-9.33625668e-12-4.83652972e+04 7.02616632e+01                   4
QMLINOOX                C  19H  33O   4     G    300.00   3500.00 1760.00      1
 6.81309948e+01 7.45379902e-02-2.47878007e-05 3.55693559e-09-1.75307126e-13    2
-8.29474454e+04-3.08878538e+02 1.76458104e-02 2.29341056e-01-1.56722232e-04    3
 5.35320989e-08-7.27405191e-12-5.89715465e+04 5.82344142e+01                   4
QMPAOOH                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.77681786e+01 6.05584838e-02-2.66377343e-05 5.63139231e-09-4.71383628e-13    2
-7.68263296e+04-1.55143375e+02 4.12866858e+00 1.35312950e-01-8.89331232e-05    3
 2.87037586e-08-3.67587894e-12-6.47161060e+04 2.69206708e+01                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   3500.00 1230.00      1
-1.30612117e+02 6.00365422e-01-4.85197519e-04 1.58690698e-07-1.80918283e-11    2
 1.24045727e+04 7.12083761e+02 2.15554530e+01 1.05511535e-01 1.18282831e-04    3
-1.68398923e-07 4.83898018e-11-2.50286496e+04-5.35376470e+01                   4
RALD3B                  C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180077e-02-2.61696720e-05 6.65382129e-09-6.35305356e-13    2
-2.14966002e+03 5.90959839e+01 7.04072885e+00-2.01204277e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381683e+00                   4
RALD3G                  C   3H   5O   1     G    300.00   3500.00 1160.00      1
-2.96412172e+00 3.83579385e-02-2.08581719e-05 5.12593560e-09-4.77571609e-13    2
 1.72028134e+03 4.58634919e+01 6.34826535e+00 6.24625900e-03 2.06655517e-05    3
-1.87382733e-08 4.66557687e-12-4.40192456e+02-4.45537170e-01                   4
RALDEST                 C   6H   9O   3     G    300.00   3500.00 1800.00      1
 1.17688624e+01 4.16586310e-02-2.02330626e-05 4.68126751e-09-4.21941087e-13    2
-4.91007178e+04-2.27507735e+01 5.76645054e+00 5.49973240e-02-3.13486401e-05    3
 8.79814806e-09-9.93730052e-13-4.69398496e+04 9.73553160e+00                   4
RBIPHENYL               C  12H   9          G    300.00   3500.00 1450.00      1
 2.67692078e+01 2.81611415e-02-6.05667723e-06-3.69378426e-10 1.67249382e-13    2
 3.92769947e+04-1.21306413e+02-1.05625108e+01 1.31145193e-01-1.12591903e-04    3
 4.86123345e-08-8.27787353e-12 5.01031931e+04 7.26686556e+01                   4
RBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1670.00      1
 1.45390319e+01 2.69797332e-02-1.09312485e-05 2.12602294e-09-1.64284673e-13    2
-3.56893368e+04-4.22613629e+01 3.26237571e+00 5.39896881e-02-3.51916871e-05    3
 1.18108288e-08-1.61410590e-12-3.19229337e+04 1.79249204e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777671e+01 3.52558917e-02-1.42493230e-05 2.76058348e-09-2.13045169e-13    2
 6.10938819e+03-7.94713741e+01-1.83523003e+00 8.26181075e-02-5.37178363e-05    3
 1.73785513e-08-2.24331848e-12 1.37820672e+04 3.58790126e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353914e-06-2.12687585e-10 1.25840459e-13    2
-3.38086418e+03-4.22339552e+01-6.42956805e+00 9.31830717e-02-9.41722601e-05    3
 5.12938173e-08-1.10712258e-11 1.12339577e+03 5.49833259e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824813e+01 2.40796407e-02-4.51347946e-06-4.25076334e-10 1.44988488e-13    2
-3.97704754e+03-4.00543783e+01-6.60757189e+00 9.15233042e-02-9.24834752e-05    3
 5.05720227e-08-1.09413374e-11 4.82664709e+02 5.62014116e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278088e+00 9.04971362e+01                   4
RDECOO                  C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
RDIPE                   C   6H  13O   1     G    300.00   3500.00 1800.00      1
 1.69549494e+01 3.45118423e-02-1.31342732e-05 2.36150213e-09-1.67133125e-13    2
-2.78147477e+04-5.54607975e+01 6.91787207e-01 7.06522027e-02-4.32512401e-05    3
 1.35159343e-08-1.71635982e-12-2.19600093e+04 3.25588287e+01                   4
RMBOOX                  C   5H   9O   4     G    300.00   3500.00 1350.00      1
 2.46557066e+01 1.60203243e-02-2.33018024e-06-2.09432791e-10 5.96256606e-14    2
-5.87318865e+04-9.28197844e+01-3.02577545e+00 9.80395304e-02-9.34626315e-05    3
 4.47942468e-08-8.27438909e-12-5.12578864e+04 4.90347050e+01                   4
RMBX                    C   5H   9O   2     G    300.00   3500.00 1800.00      1
 1.54924702e+01 2.80794103e-02-1.20573254e-05 2.49322401e-09-2.04812728e-13    2
-3.97201864e+04-5.41810445e+01 2.13573311e+00 5.77610483e-02-3.67920237e-05    3
 1.16542234e-08-1.47717375e-12-3.49117610e+04 1.81084031e+01                   4
RMCROTA                 C   5H   7O   2     G    300.00   3500.00 1430.00      1
 1.57189282e+01 1.69463336e-02-4.46708252e-06 5.66631307e-10-2.76621493e-14    2
-3.23219582e+04-4.94508733e+01 1.47581476e-01 6.05025483e-02-5.01554196e-05    3
 2.18665554e-08-3.75142509e-12-2.78685530e+04 3.12413465e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339062e+01 3.85260822e-02-1.58310821e-05 3.15191459e-09-2.53163787e-13    2
-5.89957980e+03-7.33836419e+01-9.95790329e+00 9.91745477e-02-6.63714701e-05    3
 2.18705768e-08-2.85297798e-12 3.92547162e+03 7.43253244e+01                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.27624311e+01 3.77290665e-02-1.50512076e-05 2.88934934e-09-2.22140396e-13    2
-2.53740824e+04-9.90983226e+01-6.71698823e+00 1.03238887e-01-6.96427248e-05    3
 2.31084298e-08-3.03034602e-12-1.47614915e+04 6.04504445e+01                   4
RMDOOX                  C  11H  21O   4     G    300.00   3500.00 1800.00      1
 3.96894034e+01 5.38225057e-02-2.02775001e-05 3.64793874e-09-2.61216335e-13    2
-8.38472341e+04-1.67546736e+02 4.70466765e+00 1.31566363e-01-8.50640479e-05    3
 2.76429564e-08-3.59385768e-12-7.12527292e+04 2.17979520e+01                   4
RMDX                    C  11H  21O   2     G    300.00   3500.00 1800.00      1
 2.51620868e+01 7.14154614e-02-3.28250989e-05 7.27501997e-09-6.35222696e-13    2
-5.95987259e+04-9.23572595e+01 1.85440015e+00 1.23210321e-01-7.59874815e-05    3
 2.32610876e-08-2.85550987e-12-5.12079587e+04 3.37888029e+01                   4
RME7                    C   8H  15O   2     G    300.00   3500.00 1800.00      1
 2.40410392e+01 4.26053894e-02-1.71372001e-05 3.34440554e-09-2.61909734e-13    2
-4.89929735e+04-9.20931877e+01 2.93892065e+00 8.94989861e-02-5.62151974e-05    3
 1.78177379e-08-2.27209478e-12-4.13962109e+04 2.21158799e+01                   4
RMEOLEA                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65772245e+01 8.98805970e-02-3.42288160e-05 6.24735813e-09-4.55216117e-13    2
-8.06885447e+04-2.49965378e+02-1.57106282e-01 2.15956888e-01-1.39292391e-04    3
 4.51597935e-08-5.85972103e-12-6.02641856e+04 5.70926555e+01                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   3500.00 1800.00      1
 5.68288430e+01 9.87024571e-02-3.87236246e-05 7.19531442e-09-5.31279781e-13    2
-1.23280985e+05-2.44956753e+02 2.29713937e+00 2.19884021e-01-1.39708261e-04    3
 4.45970316e-08-5.72596272e-12-1.03649572e+05 5.01802030e+01                   4
RMEOLES                 C  19H  35O   2     G    300.00   3500.00 1800.00      1
 5.65772245e+01 8.98805970e-02-3.42288160e-05 6.24735813e-09-4.55216117e-13    2
-8.06885447e+04-2.49965378e+02-1.57106282e-01 2.15956888e-01-1.39292391e-04    3
 4.51597935e-08-5.85972103e-12-6.02641856e+04 5.70926555e+01                   4
RMLIN1A                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150691e+01 7.42461115e-02-2.53824843e-05 3.82833735e-09-2.08614643e-13    2
-4.82863749e+04-2.69048825e+02-9.12524230e-01 2.08529652e-01-1.37285435e-04    3
 4.52738746e-08-5.96493926e-12-2.65324413e+04 5.79979154e+01                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   3500.00 1650.00      1
 5.48798863e+01 9.05843840e-02-3.54321193e-05 6.50176029e-09-4.69049023e-13    2
-7.13229393e+04-2.34809039e+02-1.47497564e+00 2.27202231e-01-1.59630162e-04    3
 5.66827877e-08-8.07223499e-12-5.27258349e+04 6.52917158e+01                   4
RMLIN1X                 C  19H  31O   2     G    300.00   3500.00 1800.00      1
 5.95150691e+01 7.42461115e-02-2.53824843e-05 3.82833735e-09-2.08614643e-13    2
-4.82863749e+04-2.69048825e+02-9.12524230e-01 2.08529652e-01-1.37285435e-04    3
 4.52738746e-08-5.96493926e-12-2.65324413e+04 5.79979154e+01                   4
RMLINA                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954712e+01 8.40022248e-02-3.15645422e-05 5.64019755e-09-4.00096883e-13    2
-6.69574846e+04-2.54485602e+02-1.30856133e+00 2.14011186e-01-1.39905343e-04    3
 4.57664202e-08-5.97318336e-12-4.58960329e+04 6.21504271e+01                   4
RMLINOOX                C  19H  33O   4     G    300.00   3500.00 1780.00      1
 6.32132444e+01 8.05239356e-02-2.78197745e-05 4.27200724e-09-2.39927804e-13    2
-8.77238917e+04-2.82700411e+02 1.99661323e+00 2.18089399e-01-1.43745727e-04    3
 4.76899669e-08-6.33795584e-12-6.59307710e+04 4.79327752e+01                   4
RMLINX                  C  19H  33O   2     G    300.00   3500.00 1800.00      1
 5.71954712e+01 8.40022248e-02-3.15645422e-05 5.64019755e-09-4.00096883e-13    2
-6.69574846e+04-2.54485602e+02-1.30856133e+00 2.14011186e-01-1.39905343e-04    3
 4.57664202e-08-5.97318336e-12-4.58960329e+04 6.21504271e+01                   4
RMP3                    C   4H   7O   2     G    300.00   3500.00 1800.00      1
 9.46731146e+00 2.78903391e-02-1.31079861e-05 2.94998316e-09-2.60075548e-13    2
-3.18264551e+04-1.93081295e+01 3.67472870e+00 4.07627453e-02-2.38349912e-05    3
 6.92294802e-09-8.11876222e-13-2.97411253e+04 1.20425368e+01                   4
RMPAOOX                 C  17H  33O   4     G    300.00   3500.00 1800.00      1
 3.96894034e+01 5.38225057e-02-2.02775001e-05 3.64793874e-09-2.61216335e-13    2
-8.38472341e+04-1.67546736e+02 4.70466765e+00 1.31566363e-01-8.50640479e-05    3
 2.76429564e-08-3.59385768e-12-7.12527292e+04 2.17979520e+01                   4
RMPAX                   C  17H  33O   2     G    300.00   3500.00 1570.00      1
 4.65991944e+01 8.79958559e-02-3.11818152e-05 4.72867036e-09-2.34133930e-13    2
-8.86750528e+04-2.03460488e+02-5.53001427e+00 2.20809126e-01-1.58073475e-04    3
 5.86104792e-08-8.81403979e-12-7.23064813e+04 7.15470253e+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   3500.00 1250.00      1
-1.20700825e+02 5.67736647e-01-4.52750605e-04 1.47317719e-07-1.67528750e-11    2
 1.02039730e+04 6.60024010e+02 1.91170969e+01 1.20319297e-01 8.41502162e-05    3
-1.39029386e-07 4.05165459e-11-2.47505076e+04-4.57161098e+01                   4
RMTBE                   C   5H  11O   1     G    300.00   3500.00 1370.00      1
 1.09269229e+01 3.74766266e-02-1.73062474e-05 3.86241414e-09-3.39119741e-13    2
-1.88007827e+04-2.53563680e+01-1.81069448e-01 6.99087211e-02-5.28158399e-05    3
 2.11420212e-08-3.49233271e-12-1.57571928e+04 3.17301895e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278088e+00 9.04971362e+01                   4
RSTEAX                  C  19H  37O   2     G    300.00   3500.00 1590.00      1
 5.46335802e+01 9.34230719e-02-3.19964312e-05 4.67181818e-09-2.16706943e-13    2
-9.74617261e+04-2.43777088e+02-6.34709308e+00 2.46833571e-01-1.76723317e-04    3
 6.53539506e-08-9.75792273e-12-7.80698720e+04 7.86982236e+01                   4
RTC4H8OH                C   4H   9O   1     G    300.00   3500.00 1380.00      1
 8.66823484e+00 3.01271731e-02-1.35256253e-05 2.94117291e-09-2.52822189e-13    2
-1.73478965e+04-1.68023720e+01 1.39901320e-03 5.52484364e-02-4.08313463e-05    3
 1.61323424e-08-2.64252681e-12-1.49558499e+04 2.78015457e+01                   4
RTC4H9O                 C   4H   9O   1     G    300.00   3500.00 1610.00      1
 1.16852527e+01 2.57155374e-02-1.07539562e-05 2.15924613e-09-1.71897014e-13    2
-1.72607591e+04-3.73085633e+01-2.94435988e-01 5.54787390e-02-3.84836472e-05    3
 1.36415198e-08-1.95485877e-12-1.34032994e+04 2.61916467e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835937e-02-9.17249482e-06 1.42952536e-09-8.46466186e-14    2
 3.95646504e+03-1.44540610e+02-1.09331575e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619031e+01-7.89283132e-03 1.09697206e-05-3.89489830e-09 4.38586293e-13    2
-1.76924159e+04-2.71823424e+02-1.36343924e+01 1.41210048e-01-1.13282678e-04    3
 4.21245088e-08-5.95299802e-12 6.46225047e+03 9.13157248e+01                   4
RUME10                  C  11H  19O   2     G    300.00   3500.00 1450.00      1
 2.35916369e+01 6.52041736e-02-2.68467537e-05 5.44034955e-09-4.42864735e-13    2
-3.58672705e+04-8.27430018e+01 1.64400814e+00 1.25749356e-01-8.94797013e-05    3
 3.42371070e-08-5.40782293e-12-2.95024582e+04 3.12965588e+01                   4
RUME16                  C  17H  31O   2     G    300.00   3500.00 1790.00      1
 5.62816009e+01 7.14355580e-02-2.43272135e-05 3.65699376e-09-1.98260551e-13    2
-7.53409955e+04-2.53924384e+02 9.94524607e-01 1.94982097e-01-1.27857833e-04    3
 4.22158836e-08-5.58358037e-12-5.55482222e+04 4.49927995e+01                   4
RUME7                   C   8H  13O   2     G    300.00   3500.00 1800.00      1
 1.85903431e+01 4.63199659e-02-2.12076343e-05 4.67919597e-09-4.06994657e-13    2
-3.29183962e+04-6.07637830e+01 2.66158720e+00 8.17172013e-02-5.07053305e-05    3
 1.56042686e-08-1.92436586e-12-2.71840440e+04 2.54459670e+01                   4
RXYLENE                 C   8H   9          G    300.00   3500.00 1380.00      1
 9.50606195e+00 4.15939315e-02-1.79471777e-05 3.41861978e-09-2.36020443e-13    2
 1.46969060e+04-2.59567399e+01-2.80920460e+00 7.72903563e-02-5.67476394e-05    3
 2.21628042e-08-3.63170602e-12 1.80959195e+04 3.74238465e+01                   4
SC4H7                   C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017753e+00 1.98466503e-02-6.37614062e-06 5.28652771e-10 3.81103730e-14    2
 1.19533850e+04-1.83767118e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
TAME                    C   6H  14O   1     G    300.00   3500.00 1320.00      1
 1.13309761e+01 4.74280944e-02-1.96957502e-05 3.66860750e-09-2.50688228e-13    2
-4.42745214e+04-3.17952394e+01-2.12836721e+00 8.82139832e-02-6.60433511e-05    3
 2.70764868e-08-4.68399869e-12-4.07212548e+04 3.68750527e+01                   4
TC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1440.00      1
 9.08150387e+00 3.22201837e-02-1.41979352e-05 3.03249263e-09-2.56658356e-13    2
-4.23917231e+04-2.36263218e+01-6.99999563e-01 5.93910266e-02-4.25008966e-05    3
 1.61357155e-08-2.53152343e-12-3.95746501e+04 2.71305359e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565536e-05 2.20632462e-09-1.51941206e-13    2
-9.85314330e+03-1.11161769e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576861e+01 4.50315825e-02-1.97554195e-05 4.21197817e-09-3.57314917e-13    2
-1.09025839e+04-5.35378398e+01-2.75522789e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
U2ME12                  C  13H  22O   2     G    300.00   3500.00 1610.00      1
 3.12799449e+01 7.15415882e-02-3.01181538e-05 6.08643201e-09-4.87334868e-13    2
-6.28268100e+04-1.24478592e+02 1.12650720e+00 1.46456961e-01-9.99150853e-05    3
 3.49878529e-08-4.97513315e-12-5.31174030e+04 3.53544123e+01                   4
UME10                   C  11H  20O   2     G    300.00   3500.00 1800.00      1
 3.48566736e+01 5.08631615e-02-1.90027410e-05 3.39432106e-09-2.41664061e-13    2
-7.27334602e+04-1.48477392e+02 1.08700033e+00 1.25906880e-01-8.15391729e-05    3
 2.65559625e-08-3.45855871e-12-6.05763778e+04 3.42911241e+01                   4
UME16                   C  17H  32O   2     G    300.00   3500.00 1580.00      1
 4.52339702e+01 8.65152352e-02-3.05153342e-05 4.60674378e-09-2.26752205e-13    2
-9.22046847e+04-1.94026893e+02-6.34895832e+00 2.17104928e-01-1.54492890e-04    3
 5.69179489e-08-8.50384163e-12-7.59044793e+04 7.84262324e+01                   4
UME7                    C   8H  14O   2     G    300.00   3500.00 1800.00      1
 2.58473842e+01 3.62113327e-02-1.33124030e-05 2.32937526e-09-1.61944568e-13    2
-5.91274188e+04-1.03960065e+02 2.21977808e+00 8.87171241e-02-5.70672292e-05    3
 1.85348664e-08-2.41270723e-12-5.06214805e+04 2.39174684e+01                   4
XYLENE                  C   8H  10          G    300.00   3500.00 1640.00      1
 1.72256243e+01 2.83565600e-02-6.90689954e-06-3.57091403e-10 2.09419626e-13    2
-6.87239337e+03-6.97341599e+01-5.12303971e+00 8.28654966e-02-5.67626342e-05    3
 1.99094674e-08-2.87999483e-12 4.57968429e+02 4.91410252e+01                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   3500.00 1410.00      1
 1.71509971e+01 3.21642995e-02-1.45265250e-05 3.16055984e-09-2.71089893e-13    2
-4.87167967e+04-4.94521678e+01 4.90929016e+00 6.68925461e-02-5.14714682e-05    3
 2.06286181e-08-3.36826334e-12-4.52646353e+04 1.38131161e+01                   4
ZDECA                   C  10H  17O   4     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
ZMBOOX                  C   5H   9O   6     G    300.00   3500.00 1310.00      1
 2.94016942e+01 1.57346453e-02-2.10565670e-06-2.30310175e-10 5.80528651e-14    2
-7.03637113e+04-1.09596841e+02-1.66570869e+00 1.10596944e-01-1.10726610e-04    3
 5.50475284e-08-1.04911530e-11-6.22240518e+04 4.86744607e+01                   4
ZMDOOH                  C  11H  21O   6     G    300.00   3500.00 1780.00      1
 4.89601122e+01 4.69646617e-02-1.61477773e-05 2.58757356e-09-1.58080023e-13    2
-9.96313675e+04-2.11226530e+02 6.91495056e+00 1.41448171e-01-9.57687121e-05    3
 3.24081484e-08-4.34636300e-12-8.46632899e+04 1.58608722e+01                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   3500.00 1540.00      1
 5.74950108e+01 9.92606422e-02-3.35004082e-05 5.08063679e-09-2.82240300e-13    2
-1.09648465e+05-2.38315353e+02 2.38451828e+00 2.42404779e-01-1.72926515e-04    3
 6.54382588e-08-1.00805556e-11-9.26744334e+04 5.13566583e+01                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   3500.00 1690.00      1
 6.61920071e+01 8.18444133e-02-3.03706056e-05 5.17171152e-09-3.39000627e-13    2
-8.83104294e+04-2.93138255e+02 7.95447186e-01 2.36629171e-01-1.67753526e-04    3
 5.93661575e-08-8.35593051e-12-6.62063921e+04 5.66777851e+01                   4
ZMLINOOX                C  19H  33O   6     G    300.00   3500.00 1530.00      1
 6.14087077e+01 8.58331824e-02-2.98017595e-05 4.63939709e-09-2.65661024e-13    2
-9.65914210e+04-2.81173958e+02 1.31186651e+00 2.42949107e-01-1.83836980e-04    3
 7.17571402e-08-1.12326125e-11-7.82017876e+04 3.43158089e+01                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   3500.00 1780.00      1
 4.89601122e+01 4.69646617e-02-1.61477773e-05 2.58757356e-09-1.58080023e-13    2
-9.96313675e+04-2.11226530e+02 6.91495056e+00 1.41448171e-01-9.57687121e-05    3
 3.24081484e-08-4.34636300e-12-8.46632899e+04 1.58608722e+01                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   3500.00 1250.00      1
-6.22995292e+01 3.41575945e-01-2.69706994e-04 8.71969173e-08-9.87435445e-12    2
 1.57160052e+04 3.57020399e+02 1.61954271e+01 9.03920846e-02 3.17136382e-05    3
-7.35607531e-08 2.22771796e-11-3.90773390e+03-3.91880337e+01                   4
END

