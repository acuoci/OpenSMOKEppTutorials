!***********************************************************************
!SURFACE MECHANISM FOR STEAM REFORMING AND PARTIAL OXIDATION 
!OF METHANE AND HEXADECANE OVER RHODIUM
!***********************************************************************
!****                                                                  *
!****     SR/CPO CH4/C16H34 ON RH - SURFACE MECHANISM                  *
!****                                                                  *
!****     Version 1.0, March  2008                                     *
!****     L. Maier, O. Deutschmann                                     *
!****     KIT (Karlsruhe Institute of Technology)                      *
!****     Contact: mail@detchem.com (O. Deutschmann)                   * 
!****                                                                  *
!****     References:                                                  *
!****     J. Thormann, L. Maier, P. Pfeifer, U. Kunz, K. Schubert,     *
!****     O. Deutschmann.International J. Hydrogen Energy              *
!****     34 (2009), 5108-5120                                         * 
!****     www.detchem.com/mechanisms                                   * 
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****     STICK: A in next reaction is initial sticking coefficient    *
!****                                                                  *
!****                                                                  *
!****     (SURFACE CHEMKIN format)                                     *
!****                                                                  * 
!***********************************************************************   

THERMO
   300.000  1000.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2                      N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
C16H34                  C  16H  34    0    0G   300.00   3500.00  1000.00      1
-0.82120881E+00 0.17984817E+00-0.10401813E-03 0.28694978E-07-0.29946687E-11    2
-0.51322863E+05 0.50451675E+02 0.14856790E+01 0.15814024E+00-0.25881841E-04    3
-0.73410093E-07 0.41458327E-10-0.52185547E+05 0.40077819E+02                   4
CH4               121286C   1H   4          G  0300.00   5000.00  1000.00      1
 0.01683478E+02 0.10237236E-01-0.03875128E-04 0.06785585E-08-0.04503423E-12    2
-0.10080787E+05 0.09623395E+02 0.07787415E+01 0.01747668E+00-0.02783409E-03    3
 0.03049708E-06-0.12239307E-10-0.09825229E+05 0.13722195E+02                   4
CO                121286C   1O   1          G  0300.00   5000.00  1000.00      1
 0.03025078E+02 0.14426885E-02-0.05630827E-05 0.10185813E-09-0.06910951E-13    2
-0.14268350E+05 0.06108217E+02 0.03262451E+02 0.15119409E-02-0.03881755E-04    3
 0.05581944E-07-0.02474951E-10-0.14310539E+05 0.04848897E+02                   4
CO2               121286C   1O   2          G  0300.00   5000.00  1000.00      1
 0.04453623E+02 0.03140168E-01-0.12784105E-05 0.02393996E-08-0.16690333E-13    2
-0.04896696E+06-0.09553959E+01 0.02275724E+02 0.09922072E-01-0.10409113E-04    3
 0.06866686E-07-0.02117280E-10-0.04837314E+06 0.10188488E+02                   4
H2                121286H   2               G  0300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633828E-06-0.09231578E-10 0.15827519E-14    2
-0.08350340E+04-0.13551101E+01 0.03298124E+02 0.08249441E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.10125209E+04-0.03294094E+02                   4
H2O                20387H   2O   1          G  0300.00   5000.00  1000.00      1
 0.02672145E+02 0.03056293E-01-0.08730260E-05 0.12009964E-09-0.06391618E-13    2
-0.02989921E+06 0.06862817E+02 0.03386842E+02 0.03474982E-01-0.06354696E-04    3
 0.06968581E-07-0.02506588E-10-0.03020811E+06 0.02590232E+02                   4
O2                121386O   2               G  0300.00   5000.00  1000.00      1
 0.03697578E+02 0.06135197E-02-0.12588420E-06 0.01775281E-09-0.11364354E-14    2
-0.12339301E+04 0.03189165E+02 0.03212936E+02 0.11274864E-02-0.05756150E-05    3
 0.13138773E-08-0.08768554E-11-0.10052490E+04 0.06034737E+02                   4
C_Rh                    C   1RH  1    0    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
CH_Rh                   H   1C   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00-0.00000000E+00                   4
CH2_Rh                  H   2C   1RH  1    0G   300.00    450.00   450.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E-00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E-00                   4
CH3_Rh                  H   3C   1RH  1    0G   300.00    450.00   450.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
CH4_Rh                  H   4C   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
CO_Rh                   O   1C   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
CO2_Rh                  O   2C   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
H_Rh                    H   1RH  1    0    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
H2O_Rh                  H   2O   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
HCO_Rh                  H   1O   1C   1RH  1G   300.00    450.00   450.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
O_Rh                    O   1RH  1    0    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
OH_Rh                   H   1O   1RH  1    0G   293.00   5000.00  5000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
_Rh_                    RH  1    0    0    0G   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
