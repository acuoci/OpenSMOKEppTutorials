!***********************************************************************
!SURFACE MECHANISM FOR PT-CATALYZED ABATMENT OF AUTOMOTIVE EXHAUST GASES
!***********************************************************************
!****                                                                  *
!****      C3H6/CH4/NOx/CO ON PT - SURFACE MECHANISM                   *
!****                                                                  *
!****     J. Koop, O. Deutschmann                                      *
!****     KIT (Karlsruhe Institute of Technology)                      * 
!****                                                                  *
!****     Reference:                                                   *
!****     J. Koop, O. Deutschmann                                      *  
!****     Appl. Catal.B: Environmental 91 (2009), 47-58                *
!****     Contact: mail@detchem.com (O. Deutschmann)                   * 
!****     www.detchem.com/mechanisms                                   * 
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****     STICK: A in next reaction is initial sticking coefficient    *
!****                                                                  *
!****                                                                  *
!****     (SURFACE CHEMKIN format)                                     *
!****                                                                  * 
!*********************************************************************** 

THERMO
   300.000  1000.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
C3H6                    C   3H   6    0    0G   300.00   5000.00  1000.00      1
 6.73225690E+00 1.49083360E-02-4.94989940E-06 7.21202210E-10-3.76620430E-14    2
-9.23570310E+02-1.33133480E+01 1.49330710E+00 2.09251750E-02 4.48679380E-06    3
-1.66891210E-08 7.15814650E-12 1.07482640E+03 1.61453400E+01                   4
CO                      C   1O   1    0    0G   300.00   5000.00  1000.00      1
 3.02507806E+00 1.44268852E-03-5.63082779E-07 1.01858133E-10-6.91095156E-15    2
-1.42683496E+04 6.10821772E+00 3.26245165E+00 1.51194085E-03-3.88175522E-06    3
 5.58194424E-09-2.47495123E-12-1.43105391E+04 4.84889698E+00                   4
CO2                     C   1O   2    0    0G   300.00   5000.00  1000.00      1
 4.45362282E+00 3.14016873E-03-1.27841054E-06 2.39399667E-10-1.66903319E-14    2
-4.89669609E+04-9.55395877E-01 2.27572465E+00 9.92207229E-03-1.04091132E-05    3
 6.86668678E-09-2.11728009E-12-4.83731406E+04 1.01884880E+01                   4
H2                      H   2    0    0    0G   300.00   5000.00  1000.00      1
 3.06670950E+00 5.74737550E-04 1.39383190E-08-2.54835180E-11 2.90985740E-15    2
-8.65474120E+02-1.77984240E+00 3.35535140E+00 5.01361440E-04-2.30069080E-07    3
-4.79053240E-10 4.85225850E-13-1.01916260E+03-3.54772280E+00                   4
H2O                     H   2O   1    0    0G   300.00   5000.00  1000.00      1
 2.61104720E+00 3.15631300E-03-9.29854380E-07 1.33315380E-10-7.46893510E-15    2
-2.98681670E+04 7.20912680E+00 4.16772340E+00-1.81149700E-03 5.94712880E-06    3
-4.86920210E-09 1.52919910E-12-3.02899690E+04-7.31354740E-01                   4
N2                      N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
N2O                     O   1N   2    0    0G   300.00   5000.00  1000.00      1
 4.73066790E+00 2.82582670E-03-1.15581150E-06 2.12636830E-10-1.45640870E-14    2
 8.16176820E+03-1.71510730E+00 2.61891960E+00 8.64396160E-03-6.81106240E-06    3
 2.22758770E-09-8.06503300E-14 8.75901230E+03 9.22669520E+00                   4
NO                      O   1N   1    0    0G   300.00   5000.00  1000.00      1
 3.18900000E+00 1.33822810E-03-5.28993180E-07 9.59193320E-11-6.48479320E-15    2
 9.82832900E+03 6.74581260E+00 4.04595210E+00-3.41817830E-03 7.98191900E-06    3
-6.11393160E-09 1.59190760E-12 9.74539340E+03 2.99749880E+00                   4
NO2                     O   2N   1    0    0G   300.00   5000.00  1000.00      1
 4.62407710E+00 2.52603320E-03-1.06094980E-06 1.98792390E-10-1.37993840E-14    2
 2.28999000E+03 1.33241380E+00 3.45892360E+00 2.06470640E-03 6.68660670E-06    3
-9.55567250E-09 3.61958810E-12 2.81522650E+03 8.31169830E+00                   4
O2                      O   2    0    0    0G   300.00   5000.00  1000.00      1
 3.61221390E+00 7.48531660E-04-1.98206470E-07 3.37490080E-11-2.39073740E-15    2
-1.19781510E+03 3.67033070E+00 3.78371350E+00-3.02336340E-03 9.94927510E-06    3
-9.81891010E-09 3.30318250E-12-1.06381070E+03 3.64163450E+00                   4
C_Pt                    C   1Pt  1    0    0I   300.00    900.00   900.00      1
 1.47913248E-01 1.45202051E-03 4.47050620E-06-7.41988343E-09 3.64357839E-12    2
 8.39612563E+03 4.05922946E+00 1.47913248E-01 1.45202051E-03 4.47050620E-06    3
-7.41988343E-09 3.64357839E-12 8.39612563E+03 4.05922946E+00                   4
C2H3_Pt                 C   2H   3Pt  1    0I   300.00    900.00   900.00      1
 1.00267303E+00 1.12120748E-02 1.08826725E-06-7.20229473E-09 3.28613356E-12    2
 3.80551264E+03 4.19828627E+00 1.00267303E+00 1.12120748E-02 1.08826725E-06    3
-7.20229473E-09 3.28613356E-12 3.80551264E+03 4.19828627E+00                   4
C3H4_Pt1                C   3H   4Pt  1    0I   300.00   5000.00  5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C3H5_Pt                 C   3H   5Pt  1    0I   300.00    900.00   900.00      1
 1.07734328E+00 1.86760879E-02 2.25773296E-06-1.24978251E-08 5.51492067E-12    2
-4.42512847E+02 6.78924420E+00 1.07734328E+00 1.86760879E-02 2.25773296E-06    3
-1.24978251E-08 5.51492067E-12-4.42512847E+02 6.78924420E+00                   4
C3H5_Pt1                C   3H   5Pt  1    0I   300.00    900.00   900.00      1
 4.83555099E-01 1.80358010E-02 1.05860725E-05-2.44828289E-08 1.09002865E-11    2
 8.98332516E+03 7.16225851E+00 4.83555099E-01 1.80358010E-02 1.05860725E-05    3
-2.44828289E-08 1.09002865E-11 8.98332516E+03 7.16225851E+00                   4
C3H6_Pt                 C   3H   6Pt  2    0I   300.00    900.00   900.00      1
 1.85583448E+00 2.09575461E-02-2.21362246E-06-7.09409927E-09 2.97758999E-12    2
-8.13308559E+03 4.17679549E+00 1.85583448E+00 2.09575461E-02-2.21362246E-06    3
-7.09409927E-09 2.97758999E-12-8.13308559E+03 4.17679549E+00                   4
CH_Pt                   C   1H   1Pt  1    0I   300.00    900.00   900.00      1
 3.76853374E-01 4.33007371E-03 1.26813836E-06-4.03298591E-09 1.91710002E-12    2
 1.95692528E+04 2.10382533E+00 3.76853374E-01 4.33007371E-03 1.26813836E-06    3
-4.03298591E-09 1.91710002E-12 1.95692528E+04 2.10382533E+00                   4
CH2_Pt                  C   1H   2Pt  1    0I   300.00    900.00   900.00      1
 8.33824124E-02 7.46370122E-03 1.10415461E-06-5.20153053E-09 2.18780284E-12    2
 8.36101765E+03 2.55159890E+00 8.33824124E-02 7.46370122E-03 1.10415461E-06    3
-5.20153053E-09 2.18780284E-12 8.36101765E+03 2.55159890E+00                   4
CH3_Pt                  C   1H   3Pt  1    0I   300.00    900.00   900.00      1
 8.57809745E-01 9.76143682E-03-3.41063308E-06 2.57308727E-10-3.74694697E-13    2
-4.64570142E+03 1.16541017E-01 8.57809745E-01 9.76143682E-03-3.41063308E-06    3
 2.57308727E-10-3.74694697E-13-4.64570142E+03 1.16541017E-01                   4
CH3CO_Pt                C   2H   3O   1Pt  1I   300.00    900.00   900.00      1
 2.99398937E+00 1.15976265E-02-3.66470550E-06 3.58826366E-10-4.36573914E-13    2
-2.59207895E+04-4.95181670E+00 2.99398937E+00 1.15976265E-02-3.66470550E-06    3
 3.58826366E-10-4.36573914E-13-2.59207895E+04-4.95181670E+00                   4
CO_Pt                   C   1O   1Pt  1    0I   300.00    900.00   900.00      1
 2.71277410E+00 1.59098477E-03-3.74426457E-06 5.29775390E-09-2.33787849E-12    2
-3.06782579E+04-4.40481342E+00 2.71277410E+00 1.59098477E-03-3.74426457E-06    3
 5.29775390E-09-2.33787849E-12-3.06782579E+04-4.40481342E+00                   4
CO2_Pt                  C   1O   2Pt  1    0I   300.00    900.00   900.00      1
 4.10777858E+00 2.27188590E-03-4.99101157E-06 7.57467258E-09-3.73435334E-12    2
-5.16326794E+04-9.57779283E+00 4.10777858E+00 2.27188590E-03-4.99101157E-06    3
 7.57467258E-09-3.73435334E-12-5.16326794E+04-9.57779283E+00                   4
H_Pt                    H   1Pt  1    0    0I   300.00    800.00   800.00      1
 9.90750227E-01 6.94689242E-04-2.54107153E-09-1.41451113E-10 0.00000000E+00    2
-4.51438985E+03-4.19517661E+00 9.90750227E-01 6.94689242E-04-2.54107153E-09    3
-1.41451113E-10 0.00000000E+00-4.51438985E+03-4.19517661E+00                   4
H2O_Pt                  H   2O   1Pt  1    0I   300.00    800.00   800.00      1
 3.33746420E+00 3.52784936E-04 2.42556322E-06-1.48206404E-09 0.00000000E+00    2
-3.62057980E+04-9.72027689E+00 3.33746420E+00 3.52784936E-04 2.42556322E-06    3
-1.48206404E-09 0.00000000E+00-3.62057980E+04-9.72027689E+00                   4
HCOO_Pt                 C   1H   1O   2Pt  1I   300.00    900.00   900.00      1
 2.84183375E+00 4.40992330E-03-5.96551946E-06 7.32082418E-09-3.47262183E-12    2
-1.52640070E+04-5.39553627E+00 2.84183375E+00 4.40992330E-03-5.96551946E-06    3
 7.32082418E-09-3.47262183E-12-1.52640070E+04-5.39553627E+00                   4
N_Pt                    N   1Pt  1    0    0I   300.00    900.00   900.00      1
 1.86990513E+00-3.48858712E-03 1.04315115E-05-1.15987473E-08 4.77384604E-12    2
 1.35427962E+04-1.18732173E-01 1.86990513E+00-3.48858712E-03 1.04315115E-05    3
-1.15987473E-08 4.77384604E-12 1.35427962E+04-1.18732173E-01                   4
N2O_Pt                  O   1N   2Pt  1    0I   300.00    900.00   900.00      1
 3.50833254E+00 1.39878835E-03 5.72361548E-06-8.26453214E-09 3.47126761E-12    2
 1.00055866E+04-2.79050713E+00 3.50833254E+00 1.39878835E-03 5.72361548E-06    3
-8.26453214E-09 3.47126761E-12 1.00055866E+04-2.79050713E+00                   4
NO_Pt                   O   1N   1Pt  1    0I   300.00    900.00   900.00      1
 3.02717233E+00-2.35291082E-03 7.81376243E-06-7.14290546E-09 2.24302265E-12    2
 1.37772082E+03-8.77404102E-01 3.02717233E+00-2.35291082E-03 7.81376243E-06    3
-7.14290546E-09 2.24302265E-12 1.37772082E+03-8.77404102E-01                   4
NO2_Pt                  O   2N   1Pt  1    0I   300.00    900.00   900.00      1
 3.95654168E+00-8.30664675E-04 6.68591838E-06-6.06096773E-09 1.53311776E-12    2
-1.07963532E+03 5.56565050E-01 3.95654168E+00-8.30664675E-04 6.68591838E-06    3
-6.06096773E-09 1.53311776E-12-1.07963532E+03 5.56565050E-01                   4
O_Pt                    O   1Pt  1    0    0I   300.00    800.00   800.00      1
 1.52967014E+00-2.63766497E-04 1.28966071E-06-8.04441298E-10 0.00000000E+00    2
-1.40432598E+04-3.37596736E+00 1.52967014E+00-2.63766497E-04 1.28966071E-06    3
-8.04441298E-10 0.00000000E+00-1.40432598E+04-3.37596736E+00                   4
OH_Pt                   H   1O   1Pt  1    0I   300.00    800.00   800.00      1
 2.33488520E+00 3.22820417E-04 1.77158426E-06-1.19563622E-09 0.00000000E+00    2
-2.57097938E+04-7.40908407E+00 2.33488520E+00 3.22820417E-04 1.77158426E-06    3
-1.19563622E-09 0.00000000E+00-2.57097938E+04-7.40908407E+00                   4
_Pt_                    Pt  1    0    0    0I   300.00   5000.00  5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
