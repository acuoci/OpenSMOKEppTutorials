!*********************************************************************
!SURFACE MECHANISM OF THE C2H6-O2 REACTION ON PT                     *
!*********************************************************************
!****                                                                *
!****     C2H6 - O2 SURFACE MECHANISM ON PT                          *
!****                                                                *
!****     D. Zerkle, Los Alamos National Laboratory, USA             *
!****     O. Deutschmann, M. Wolf, Heidelberg University, Germany    *
!****                                                                *
!****     Ref.: D.K. Zerkle, M.D. Allendorf, M. Wolf, O. Deutschmann.*
!****           Understanding Homogeneous and Heterogeneous          *
!****           Contributions to the Platinum-Catalyzed Partial      *
!****           Oxidation of Ethane in a Short Contact Time Reactor. *
!****           J. Catal. 196(2000) 18-39.                           *  
!****           (NOTE: Typos for A of Rxns 26,29,57,59 in Ref.)      *
!****                                                                *
!****     Contact: mail@detchem.com (O. Deutschmann)                 *
!****                                                                *
!****                                                                *
!****     Kinetic data:                                              *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea *
!****                                       (cm,mol,s)    -    J/mol *
!****                                                                *
!****     STICK: A in next reaction is initial sticking coefficient  *
!****                                                                *
!****     $..  : additional coverage dependence of Ea (3rd column)   *
!****               or changed reaction order (2nd column)           *
!****                                                                *
!****      see manuals on www.detchem.com for details                *
!****                                                                *
!****                                                                *
!****     Surface site density: 2.72E-9 mol/cm**2                    *
!****                                                                *
!****                                                                *
!****     CHEMKIN format Februar 2006, tested with Version 4.0.1     *
!****     Ref.: http://www.detchem.com                               *
!****                                                                *
!****                                                                *
!*********************************************************************

THERMO
   300.000  1000.000  3000.000

H2                121286H   2               G   300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633828E-06-0.09231578E-10 0.15827519E-14    2
-0.08350340E+04-0.13551101E+01 0.03298124E+02 0.08249441E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.10125209E+04-0.03294094E+02                   4
H                 120186H   1               G  0300.00   5000.00  1000.00      1
 0.02500000E+02 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.02547162E+06-0.04601176E+01 0.02500000E+02 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.02547162E+06-0.04601176E+01                   4
CH4               121286C   1H   4          G  0300.00   5000.00  1000.00      1
 0.01683478E+02 0.10237236E-01-0.03875128E-04 0.06785585E-08-0.04503423E-12    2
-0.10080787E+05 0.09623395E+02 0.07787415E+01 0.01747668E+00-0.02783409E-03    3
 0.03049708E-06-0.12239307E-10-0.09825229E+05 0.13722195E+02                   4
CH3               121286C   1H   3          G  0300.00   5000.00  1000.00      1
 0.02844051E+02 0.06137974E-01-0.02230345E-04 0.03785161E-08-0.02452159E-12    2
 0.16437809E+05 0.05452697E+02 0.02430442E+02 0.11124099E-01-0.01680220E-03    3
 0.16218288E-07-0.05864952E-10 0.16423781E+05 0.06789794E+02                   4
CHO      HCO      121286H   1C   1O   1     G  0300.00   5000.00  1000.00      1
 0.03557271E+02 0.03345572E-01-0.13350060E-05 0.02470572E-08-0.01713850E-12    2
 0.03916324E+05 0.05552299E+02 0.02898329E+02 0.06199146E-01-0.09623084E-04    3
 0.10898249E-07-0.04574885E-10 0.04159922E+05 0.08983614E+02                   4
CH2O              121286C   1H   2O   1     G  0300.00   5000.00  1000.00      1
 0.02995606E+02 0.06681321E-01-0.02628954E-04 0.04737153E-08-0.03212517E-12    2
-0.15320369E+05 0.06912572E+02 0.16527311E+01 0.12631439E-01-0.01888168E-03    3
 0.02050031E-06-0.08413237E-10-0.14865404E+05 0.13784820E+02                   4
CO2               121286C   1O   2          G  0300.00   5000.00  1000.00      1
 0.04453623E+02 0.03140168E-01-0.12784105E-05 0.02393996E-08-0.16690333E-13    2
-0.04896696E+06-0.09553959E+01 0.02275724E+02 0.09922072E-01-0.10409113E-04    3
 0.06866686E-07-0.02117280E-10-0.04837314E+06 0.10188488E+02                   4
CO                121286C   1O   1          G  0300.00   5000.00  1000.00      1
 0.03025078E+02 0.14426885E-02-0.05630827E-05 0.10185813E-09-0.06910951E-13    2
-0.14268350E+05 0.06108217E+02 0.03262451E+02 0.15119409E-02-0.03881755E-04    3
 0.05581944E-07-0.02474951E-10-0.14310539E+05 0.04848897E+02                   4
O2                121386O   2               G  0300.00   5000.00  1000.00      1
 0.03697578E+02 0.06135197E-02-0.12588420E-06 0.01775281E-09-0.11364354E-14    2
-0.12339301E+04 0.03189165E+02 0.03212936E+02 0.11274864E-02-0.05756150E-05    3
 0.13138773E-08-0.08768554E-11-0.10052490E+04 0.06034737E+02                   4
O                 120186O   1               G  0300.00   5000.00  1000.00      1
 0.02542059E+02-0.02755061E-03-0.03102803E-07 0.04551067E-10-0.04368051E-14    2
 0.02923080E+06 0.04920308E+02 0.02946428E+02-0.16381665E-02 0.02421031E-04    3
-0.16028431E-08 0.03890696E-11 0.02914764E+06 0.02963995E+02                   4
OH                121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 0.03886888E+05 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 0.03606781E+05 0.13588605E+01                   4
HO2                20387H   1O   2          G  0300.00   5000.00  1000.00      1
 0.04072191E+02 0.02131296E-01-0.05308145E-05 0.06112269E-09-0.02841164E-13    2
-0.15797270E+03 0.03476029E+02 0.02979963E+02 0.04996697E-01-0.03790997E-04    3
 0.02354192E-07-0.08089024E-11 0.01762273E+04 0.09222724E+02                   4
H2O2              120186H   2O   2          G  0300.00   5000.00  1000.00      1
 0.04573167E+02 0.04336136E-01-0.14746888E-05 0.02348903E-08-0.14316536E-13    2
-0.01800696E+06 0.05011369E+01 0.03388753E+02 0.06569226E-01-0.14850125E-06    3
-0.04625805E-07 0.02471514E-10-0.01766314E+06 0.06785363E+02                   4
H2O                20387H   2O   1          G  0300.00   5000.00  1000.00      1
 0.02672145E+02 0.03056293E-01-0.08730260E-05 0.12009964E-09-0.06391618E-13    2
-0.02989921E+06 0.06862817E+02 0.03386842E+02 0.03474982E-01-0.06354696E-04    3
 0.06968581E-07-0.02506588E-10-0.03020811E+06 0.02590232E+02                   4
C2H2              121386C   2H   2          G  0300.00   5000.00  1000.00      1
 0.04436770E+02 0.05376039E-01-0.01912816E-04 0.03286379E-08-0.02156709E-12    2
 0.02566766E+06-0.02800338E+02 0.02013562E+02 0.15190446E-01-0.16163189E-04    3
 0.09078992E-07-0.01912746E-10 0.02612444E+06 0.08805378E+02                   4
C2H3               12787C   2H   3          G  0300.00   5000.00  1000.00      1
 0.05933468E+02 0.04017745E-01-0.03966739E-05-0.14412666E-09 0.02378643E-12    2
 0.03185434E+06-0.08530313E+02 0.02459276E+02 0.07371476E-01 0.02109872E-04    3
-0.13216421E-08-0.11847838E-11 0.03335225E+06 0.11556202E+02                   4
C2H4              121286C   2H   4          G  0300.00   5000.00  1000.00      1
 0.03528418E+02 0.11485185E-01-0.04418385E-04 0.07844600E-08-0.05266848E-12    2
 0.04428288E+05 0.02230389E+02-0.08614880E+01 0.02796162E+00-0.03388677E-03    3
 0.02785152E-06-0.09737879E-10 0.05573046E+05 0.02421148E+03                   4
C2H5               12387C   2H   5          G  0300.00   5000.00  1000.00      1
 0.07190480E+02 0.06484077E-01-0.06428064E-05-0.02347879E-08 0.03880877E-12    2
 0.10674549E+05-0.14780892E+02 0.02690701E+02 0.08719133E-01 0.04419838E-04    3
 0.09338703E-08-0.03927773E-10 0.12870404E+05 0.12138195E+02                   4
C2H6              121686C   2H   6          G  0300.00   4000.00  1000.00      1
 0.04825938E+02 0.13840429E-01-0.04557258E-04 0.06724967E-08-0.03598161E-12    2
-0.12717793E+05-0.05239506E+02 0.14625388E+01 0.15494667E-01 0.05780507E-04    3
-0.12578319E-07 0.04586267E-10-0.11239176E+05 0.14432295E+02                   4
CH2CO             121686C   2H   2O   1     G  0300.00   5000.00  1000.00      1
 0.06038817E+02 0.05804840E-01-0.01920953E-04 0.02794484E-08-0.14588676E-13    2
-0.08583402E+05-0.07657581E+02 0.02974970E+02 0.12118712E-01-0.02345045E-04    3
-0.06466685E-07 0.03905649E-10-0.07632636E+05 0.08673553E+02                   4
CH2CHO  OH3C2     T04/83O   1H   3C   2    0G   300.     5000.    1000.00     R1
 0.59756699E+01 0.81305914E-02-0.27436245E-05 0.40703041E-09-0.21760171E-13    2
 0.49032178E+03-0.50452509E+01 0.34090624E+01 0.10738574E-01 0.18914925E-05    3
 0.71585831E-08 0.28673851E-11 0.15214766E+04 0.95582905E+01           1552.7  4
CH3O              121686C   1H   3O   1     G  0300.00   3000.00  1000.00      1
 0.03770799E+02 0.07871497E-01-0.02656384E-04 0.03944431E-08-0.02112616E-12    2
 0.12783252E+03 0.02929575E+02 0.02106204E+02 0.07216595E-01 0.05338472E-04    3
-0.07377636E-07 0.02075610E-10 0.09786011E+04 0.13152177E+02                   4
CH2      CH2      120186C   1H   2          G  0250.00   4000.00  1000.00      1
 0.03636407E+02 0.01933056E-01-0.01687016E-05-0.10098994E-09 0.01808255E-12    2
 0.04534134E+06 0.02156560E+02 0.03762237E+02 0.11598191E-02 0.02489585E-05    3
 0.08800836E-08-0.07332435E-11 0.04536790E+06 0.01712577E+02                   4
HCCO               32387H   1C   2O   1     G  0300.00   4000.00  1000.00      1
 0.06758073E+02 0.02000400E-01-0.02027607E-05-0.10411318E-09 0.01965164E-12    2
 0.01901513E+06-0.09071262E+02 0.05047965E+02 0.04453478E-01 0.02268282E-05    3
-0.14820945E-08 0.02250741E-11 0.01965891E+06 0.04818439E+01                   4
N2                121286N   2               G  0300.00   5000.00  1000.00      1
 0.02926640E+02 0.14879768E-02-0.05684760E-05 0.10097038E-09-0.06753351E-13    2
-0.09227977E+04 0.05980528E+02 0.03298677E+02 0.14082404E-02-0.03963222E-04    3
 0.05641515E-07-0.02444854E-10-0.10208999E+04 0.03950372E+02                   4
_Pt_       dummy        PT  1               S   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H_Pt                   0H   1PT  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
O_Pt                   0O   1PT  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
OH_Pt                  0O   1H   1PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O_Pt                 0O   1H   2PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C_Pt                   0C   1PT  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO_Pt       dummy      0C   1O   1PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO2_Pt      dummy      0C   1O   2PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH3_Pt                 0C   1H   3PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH2_Pt                 0C   1H   2PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH_Pt                  0C   1H   1PT  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H6_Pt2               0C   2H   6PT  2     I   300.0    3000.0   1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H5_Pt                0C   2H   5PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H4_Pt2               0C   2H   4PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H4_Pt1               0C   2H   4PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H3_Pt2               0C   2H   3PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H3_Pt1               0C   2H   3PT  1     I   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H2_Pt3               0C   2H   2PT  1     I   300.0    3000.0   1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H2_Pt1               0C   2H   2PT  1     I   300.0    3000.0   1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H_Pt1                0C   2H   1PT  1     I   300.0    3000.0   1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
