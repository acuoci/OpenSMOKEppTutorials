!***********************************************************************
!SURFACE MECHANISM FOR STEAM REFORMING AND PARTIAL OXIDATION OF METHANE 
!OVER RHODIUM
!***********************************************************************
!****                                                                  *
!****     SR/CPO CH4 ON RH - SURFACE MECHANISM                         *
!****                                                                  *
!****     Version 2.0, March  2008                                     *
!****     L. Maier, O. Deutschmann                                     *
!****     KIT (Karlsruhe Institute of Technology)                      *
!****     Contact: mail@detchem.com (O. Deutschmann)                   * 
!****                                                                  *
!****     References:                                                  *
!****     J. Thormann, L. Maier, P. Pfeifer, U. Kunz, K. Schubert,     *
!****     O. Deutschmann.International J. Hydrogen Energy              *
!****     34 (2009), 5108-5120                                         * 
!****     www.detchem.com/mechanisms                                   * 
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****     STICK: A in next reaction is initial sticking coefficient    *
!****                                                                  *
!****                                                                  *
!****     (SURFACE CHEMKIN format)                                     *
!****                                                                  * 
!*********************************************************************** 

THERMO
   300.000  1000.000  3000.000

CH4                     C   1H   4    0     G   300.00   5000.00  1000.00      1
 0.16834780E+01 0.10237236E-01-0.38751280E-05 0.67855850E-09-0.45034230E-13    2
-0.10080787E+05 0.96233950E+01 0.77874150E+00 0.17476680E-01-0.27834090E-04    3
 0.30497080E-07-0.12239307E-10-0.98252290E+04 0.13722195E+02                   4
O2                      O   2    0    0     G   300.00   5000.00  1000.00      1
 0.36975780E+01 0.61351970E-03-0.12588420E-06 0.17752810E-10-0.11364354E-14    2
-0.12339301E+04 0.31891650E+01 0.32129360E+01 0.11274864E-02-0.57561500E-06    3
 0.13138773E-08-0.87685540E-12-0.10052490E+04 0.60347370E+01                   4
CO                      C   1O   1    0     G   300.00   5000.00  1000.00      1
 0.30250780E+01 0.14426885E-02-0.56308270E-06 0.10185813E-09-0.69109510E-14    2
-0.14268350E+05 0.61082170E+01 0.32624510E+01 0.15119409E-02-0.38817550E-05    3
 0.55819440E-08-0.24749510E-11-0.14310539E+05 0.48488970E+01                   4
CO2                     C   1O   2    0     G   300.00   5000.00  1000.00      1
 0.44536230E+01 0.31401680E-02-0.12784105E-05 0.23939960E-09-0.16690333E-13    2
-0.48966960E+05-0.95539590E+00 0.22757240E+01 0.99220720E-02-0.10409113E-04    3
 0.68666860E-08-0.21172800E-11-0.48373140E+05 0.10188488E+02                   4
H2                      H   2    0    0     G   300.00   5000.00  1000.00      1
 0.29914230E+01 0.70006440E-03-0.56338280E-07-0.92315780E-11 0.15827519E-14    2
-0.83503400E+03-0.13551101E+01 0.32981240E+01 0.82494410E-03-0.81430150E-06    3
-0.94754340E-10 0.41348720E-12-0.10125209E+04-0.32940940E+01                   4
H2O                     H   2O   1    0     G   300.00   5000.00  1000.00      1
 0.26721450E+01 0.30562930E-02-0.87302600E-06 0.12009964E-09-0.63916180E-14    2
-0.29899210E+05 0.68628170E+01 0.33868420E+01 0.34749820E-02-0.63546960E-05    3
 0.69685810E-08-0.25065880E-11-0.30208110E+05 0.25902320E+01                   4
N2                      N   2    0    0     G   300.00   5000.00  1000.00      1
 0.29266400E+01 0.14879768E-02-0.56847600E-06 0.10097038E-09-0.67533510E-14    2
-0.92279770E+03 0.59805280E+01 0.32986770E+01 0.14082404E-02-0.39632220E-05    3
 0.56415150E-08-0.24448540E-11-0.10208999E+04 0.39503720E+01                   4
 
RH(s)                   RH  1    0    0     G   300.00   3000.00  1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O(s)                  H   2O   1RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
H(s)                    H   1RH  1    0     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
OH(s)                   H   1O   1RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(s)                   C   1O   1RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
C(s)                    C   1RH  1    0     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
CH3(s)                  C   1H   3RH  1     G   300.00    450.00   450.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
CH2(s)                  C   1H   2RH  1     G   300.00    450.00   450.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
CH(s)                   C   1H   1RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00-0.00000000E+00                   4
CH4(s)                  C   1H   4RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
O(s)                    O   1RH  1    0     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
CO2(s)                  C   1O   2RH  1     G   293.00   5000.00  5000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4
HCO(s)                  C   1H   1O   1RH  1G   300.00    450.00  450.00       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00 0.00000000E+00                   4

END
