!***********************************************************************
!SURFACE MECHANISM FOR PARTIAL OXIDATION/REFORMING OF PROPANE AND 
!ISOOCTANE OVER RHODIUM
!***********************************************************************
!****                                                                  *
!****     CPO C3H8/isoC8H18 ON RH - SURFACE MECHANISM                  *
!****                                                                  *
!****     Version 1.0, Januar  2010                                    *
!****     L. Maier, M. Hartmann, O. Deutschmann                        *
!****     KIT (Karlsruhe Institute of Technology)                      *
!****     Contact: mail@detchem.com (O. Deutschmann)                   * 
!****                                                                  *
!****     References:                                                  *
!****     M. Hartmann, L. Maier, O. Deutschmann                        * 
!****     Combustion and Flame, 157 (2010) 1771-1782.                  *  
!****     www.detchem.com/mechanisms                                   * 
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****     STICK: A in next reaction is initial sticking coefficient    *
!****                                                                  *
!****                                                                  *
!****     (SURFACE CHEMKIN format)                                     *
!****                                                                  * 
!*********************************************************************** 

THERMO
   300.000  1000.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2                      N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
C3H8              120186C   3H   8          G  0300.00   5000.00  1000.00      1
 0.07525217E+02 0.01889034E+00-0.06283924E-04 0.09179373E-08-0.04812410E-12    2
-0.01646455E+06-0.01784390E+03 0.08969208E+01 0.02668986E+00 0.05431425E-04    3
-0.02126001E-06 0.09243330E-10-0.01395492E+06 0.01935533E+03                   4
CH4               121286C   1H   4          G  0300.00   5000.00  1000.00      1
 0.01683479E+02 0.01023724E+00-0.03875129E-04 0.06785585E-08-0.04503423E-12    2
-0.01008079E+06 0.09623395E+02 0.07787415E+01 0.01747668E+00-0.02783409E-03    3
 0.03049708E-06-0.01223931E-09-0.09825229E+05 0.01372219E+03                   4
CO                121286C   1O   1          G  0300.00   5000.00  1000.00      1
 0.03025078E+02 0.01442689E-01-0.05630828E-05 0.01018581E-08-0.06910952E-13    2
-0.01426835E+06 0.06108218E+02 0.03262452E+02 0.01511941E-01-0.03881755E-04    3
 0.05581944E-07-0.02474951E-10-0.01431054E+06 0.04848897E+02                   4
CO2               121286C   1O   2          G  0300.00   5000.00  1000.00      1
 0.04453623E+02 0.03140169E-01-0.01278411E-04 0.02393997E-08-0.01669033E-12    2
-0.04896696E+06-0.09553959E+01 0.02275725E+02 0.09922072E-01-0.01040911E-03    3
 0.06866687E-07-0.02117280E-10-0.04837314E+06 0.01018849E+03                   4
H2                121286H   2               G  0300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633829E-06-0.09231578E-10 0.01582752E-13    2
-0.08350340E+04-0.01355110E+02 0.03298124E+02 0.08249442E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.01012521E+05-0.03294094E+02                   4
H2O                20387H   2O   1          G  0300.00   5000.00  1000.00      1
 0.02672146E+02 0.03056293E-01-0.08730260E-05 0.01200996E-08-0.06391618E-13    2
-0.02989921E+06 0.06862817E+02 0.03386842E+02 0.03474982E-01-0.06354696E-04    3
 0.06968581E-07-0.02506588E-10-0.03020811E+06 0.02590233E+02                   4
I-C8H18     RANZI       C   8H  18          G  0300.00   5000.00  1388.00      1
  .17556581E+02 0.49924288E-01 -.17202017E-04  .27551890E-08 -.16941933E-12    2
 -.36369008E+05 -.67112610E+02 -.20321865E+01  .94684526E-01 -.35743305E-04    3
 -.16594676E-07  .12534632E-10 -.30683273E+05  .35986145E+02                   4
O2                121386O   2               G  0300.00   5000.00  1000.00      1
 0.03697578E+02 0.06135197E-02-0.01258842E-05 0.01775281E-09-0.01136435E-13    2
-0.01233930E+05 0.03189166E+02 0.03212936E+02 0.01127486E-01-0.05756150E-05    3
 0.01313877E-07-0.08768554E-11-0.01005249E+05 0.06034738E+02                   4
C_Rh                   0C   1Rh  1          S    300.00   3000.00 1000.00      1
 0.15792824E+01 0.36528701E-03-0.50657672E-07-0.34884855E-10 0.88089699E-14    2
 0.99535752E+04-0.30240495E+01 0.58924019E+00 0.25012842E-02-0.34229498E-06    3
-0.18994346E-08 0.10190406E-11 0.10236923E+05 0.21937017E+01                   4
C2H3_Rh                0C   2H   3Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
C3H6_Rh                0C   3H   6Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
C3H7_Rh                0C   3H   7Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
C3H8_Rh                0C   3H   8Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
CH_Rh                  0C   1H   1Rh  1     S    300.00   3000.00 1000.00      1
-0.48242472E-02 0.30446239E-02-0.16066099E-06-0.29041700E-09 0.57999924E-13    2
 0.22595219E+05 0.56677818E+01 0.84157485E+00 0.13095380E-02 0.28464575E-06    3
 0.63862904E-09-0.42766658E-12 0.22332801E+05 0.11452305E+01                   4
CH2_Rh                 0C   1H   2Rh  1     S    300.00   3000.00 1000.00      1
 0.74076122E+00 0.48032533E-02-0.32825633E-06-0.47779786E-09 0.10073452E-12    2
 0.10443752E+05 0.40842086E+00-0.14876404E+00 0.51396289E-02 0.11211075E-05    3
-0.82755452E-09-0.44572345E-12 0.10878700E+05 0.57451882E+01                   4
CH3_Rh                 0C   1H   3Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
CH4_Rh                 0C   1H   4Rh  1     S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
CO_Rh                  0C   1O   1Rh  1     S    300.00   3000.00 1000.00      1
 0.47083778E+01 0.96037297E-03-0.11805279E-06-0.76883826E-10 0.18232000E-13    2
-0.32311723E+05-0.16719593E+02 0.48907466E+01 0.68134235E-04 0.19768814E-06    3
 0.12388669E-08-0.90339249E-12-0.32297836E+05-0.17453161E+02                   4
CO2_Rh            081292C   1O   2Rh  1     S   300.00   3000.00  1000.00      1
 0.46900000E+00 0.62660000E-02 0.00000000E-00 0.00000000E-00 0.00000000E-00    2
-0.50458700E+05-0.45550000E+01 0.46900000E+00 0.62662000E-02 0.00000000E-00    3
 0.00000000E-00 0.00000000E-00-0.50458700E+05-0.45550000E+01                   4
H_Rh               92491H   1Rh  1          I    300.00   3000.00 1000.00      1
 0.10696996E+01 0.15432230E-02-0.15500922E-06-0.16573165E-09 0.38359347E-13    2
-0.50546128E+04-0.71555238E+01-0.13029877E+01 0.54173199E-02 0.31277972E-06    3
-0.32328533E-08 0.11362820E-11-0.42277075E+04 0.58743238E+01                   4
H2O_Rh             92491O   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.25803051E+01 0.49570827E-02-0.46894056E-06-0.52633137E-09 0.11998322E-12    2
-0.38302234E+05-0.17406322E+02-0.27651553E+01 0.13315115E-01 0.10127695E-05    3
-0.71820083E-08 0.22813776E-11-0.36398055E+05 0.12098145E+02                   4
HCO_Rh                  C   1H   1O   1Rh  1S    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
O_Rh               92491O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.19454180E+01 0.91761647E-03-0.11226719E-06-0.99099624E-10 0.24307699E-13    2
-0.14005187E+05-0.11531663E+02-0.94986904E+00 0.74042305E-02-0.10451424E-05    3
-0.61120420E-08 0.33787992E-11-0.13209912E+05 0.36137905E+01                   4
OH_Rh              92491O   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.18249973E+01 0.32501565E-02-0.31197541E-06-0.34603206E-09 0.79171472E-13    2
-0.26685492E+05-0.12280891E+02-0.20340881E+01 0.93662683E-02 0.66275214E-06    3
-0.52074887E-08 0.17088735E-11-0.25319949E+05 0.89863186E+01                   4
_Rh_                    Rh  1               S    300.0    3000.0  1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
