THERMO ALL
270.   1000.   3500. 
! NEW PHENYLACETYLENE
C6H5CCC6H5       CBS-QB3C  14H  10    0    0G   300.000  5000.000 1400.00      1 !FROM HAMADI 2022
 3.24080059E+01 3.15223030E-02-1.08906881E-05 1.70278712E-09-9.92957496E-14    2
 3.46385999E+04-1.49912722E+02-9.02216348E+00 1.40229425E-01-1.21743881E-04    3
 5.34760686E-08-9.35416414E-12 4.77334990E+04 6.81960895E+01                   4
C13H8CH2         CBS-QB3C  14H  10    0    0G   300.000  5000.000 1400.00      1 !FROM HAMADI 2022
 3.28469542E+01 3.16630850E-02-1.09601031E-05 1.71588858E-09-1.00153304E-13    2
 1.69163469E+04-1.57867490E+02-1.10527644E+01 1.47504519E-01-1.29658655E-04    3
 5.73541044E-08-1.00702016E-11 3.07102768E+04 7.29834464E+01                   4
C5H6OH                  C   5H   7O   1     G     200.0    3000.0  1000.0      1 !LPM AUTOMECH- CCSD(T)/CBS//B2PLYPD3/6-311+G(D,P) W1 IN QIAN PES, NOT MOST STABLE (W24 IS)
 7.44306564E+00 3.19941916E-02-1.57395020E-05 3.77115170E-09-3.56263749E-13    2
-3.43765939E+03-1.25591310E+01 3.45077169E+00 1.80063881E-02 6.60589621E-05    3
-1.05621589E-07 4.52181108E-11-1.48430801E+03 1.31778834E+01                   4
AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013931e+00-3.98290200e-07 3.45886082e-10-1.18293971e-13 1.38553174e-17    2
-7.45407891e+02 4.37897362e+00 2.49974489e+00 1.52569132e-06-3.17359231e-09    3
 2.74307057e-12-8.58511922e-16-7.45343207e+02 4.38079817e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811579e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324662e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42576298e-07 4.63926302e-10-1.57302170e-13 1.82971406e-17    2
-7.45426807e+02 9.27648988e-01 2.49964853e+00 2.08151569e-06-4.16682427e-09    3
 3.47465907e-12-1.04992675e-15-7.45332012e+02 9.30248556e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873259e-03 1.24226233e-06-4.19011898e-10 4.75543793e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529274e-03-1.27163634e-05    3
 1.28749173e-08-4.70027749e-12-9.43236614e+02-5.12231102e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406828e-07 6.39345346e-10-2.12551791e-13 2.44479191e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164046e-06-5.92759759e-09    3
 4.87810165e-12-1.45539320e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556201e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740147e-03 9.80122558e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959644e-04 1.33918546e-07-3.85875896e-11 4.38918689e-15    2
 2.92061519e+04 4.48358519e+00 3.14799201e+00-3.11174065e-03 6.18137897e-06    3
-5.63808798e-09 1.94866016e-12 2.91309118e+04 2.13446549e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218862e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710799e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805705e-03 5.06678941e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255381e+00 1.87486886e-03-8.59711926e-07 1.91200070e-10-1.67855286e-14    2
-1.41723335e+04 7.41443560e+00 3.75723891e+00-2.14465241e-03 5.42079005e-06    3
-4.17025963e-09 1.11901127e-12-1.43575530e+04 2.79976799e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876468e+00 2.62914704e-03-9.30606462e-07 1.43892920e-10-7.62581414e-15    2
-4.90562639e+04-2.34976452e+00 2.31684347e+00 9.22755036e-03-7.75654093e-06    3
 3.28225360e-09-5.48722482e-13-4.83626067e+04 1.00786234e+01                   4
HOCO                    H   1C   1O   2     G    200.00   3500.00 1570.00      1
 5.88810541e+00 3.28985507e-03-9.88703861e-07 1.12295277e-10-2.32818718e-15    2
-2.40914384e+04-5.05613727e+00 2.36661498e+00 1.22618052e-02-9.56063074e-06    3
 3.75217930e-09-5.81927554e-13-2.29856904e+04 1.35214769e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346405e-01 1.23697845e-02-4.99807922e-06 1.04392765e-09-8.62897416e-14    2
-9.58982501e+03 1.61752775e+01 5.23967335e+00-1.46835123e-02 5.29732711e-05    3
-5.41668822e-08 1.96318566e-11-1.02526308e+04-4.97649748e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805104e+00 6.15233477e-03-2.21179349e-06 3.74402648e-10-2.48151349e-14    2
 1.65862829e+04 5.77899818e+00 3.47829310e+00 3.54764773e-03 1.47408440e-06    3
-1.94375955e-09 5.21921232e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272972e+00 3.55431388e-03-1.28768523e-06 2.21273744e-10-1.48738147e-14    2
 4.62073492e+04 6.64284652e+00 3.76489460e+00 1.43839191e-03 4.75583077e-07    3
-4.31788591e-10 7.58292874e-14 4.58645699e+04 1.48953153e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468307e-03-1.35589914e-06 2.74980411e-10-2.36795472e-14    2
 5.06429079e+04 6.11646383e+00 4.18185434e+00-2.21134314e-03 7.71527541e-06    3
-5.95950381e-09 1.58314628e-12 5.03669407e+04-7.03002602e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472531e+00 3.92839476e-05-6.70014980e-08 3.71818694e-11-5.07306885e-15    2
 8.54504422e+04 4.79314254e+00 2.54495192e+00-2.47725281e-04 5.48018277e-07    3
-5.48551250e-10 2.04117331e-13 8.54434105e+04 4.56874273e+00                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990128e+00 2.16985238e-03-7.07637885e-07 1.23973494e-10-9.56348515e-15    2
 7.11059412e+04 8.77326061e+00 3.77264332e+00-1.58547350e-03 2.83512238e-06    3
-1.36146058e-09 2.23995332e-13 7.06312492e+04 8.79407904e-01                   4
CH3O2H                  C   1H   4O   2     G    300.00   3500.00 1090.00      1
 7.33435519e+00 9.33238534e-03-3.40995713e-06 5.79327692e-10-3.79241109e-14    2
-1.81046374e+04-1.19553974e+01 7.70006797e-01 3.34217373e-02-3.65604414e-05    3
 2.08548532e-08-4.68827401e-12-1.66736094e+04 2.02794895e+01                   4
CH3O2                   C   1H   3O   2     G    300.00   3500.00 1800.00      1
 5.64141817e+00 8.74328281e-03-3.21961406e-06 5.43695218e-10-3.45015008e-14    2
-1.19010148e+03-3.41914683e+00 1.44289632e+00 1.80733314e-02-1.09946545e-05    3
 3.42333984e-09-4.34452142e-13 3.21366390e+02 1.93041293e+01                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701530e+00 1.21538353e-02-5.02107031e-06 1.01068070e-09-8.18460823e-14    2
-2.57693409e+04 9.47420540e+00 8.47330479e-01 1.63086904e-02-8.48344961e-06    3
 2.29304341e-09-2.59952013e-13-2.50962544e+04 1.95933297e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238062e+00 5.90227637e-03-1.80340720e-06 2.13335009e-10-5.61816409e-15    2
-7.86252225e+01-7.49173677e+00 8.89660985e-01 1.70119767e-02-1.13807351e-05    3
 3.88280928e-09-5.32841479e-13 1.60316121e+03 1.85001134e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534950e+00 6.02727059e-03-2.11386821e-06 3.36085905e-10-2.00987482e-14    2
-4.03584143e+03-1.57524073e+00 2.34821579e+00 1.39600168e-02-1.08632206e-05    3
 4.62498416e-09-8.08499162e-13-3.30222106e+03 1.22661977e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335652e+00 1.00905183e-02-5.12952562e-06 1.25425207e-09-1.19639109e-13    2
-1.39080170e+04 1.59916144e+01 4.32621296e+00-7.01151853e-03 3.15176961e-05    3
-3.36478638e-08 1.23454023e-11-1.43270169e+04 2.62028902e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278258e-03-2.69184211e-06 7.21357798e-10-7.43521409e-14    2
 4.05725330e+03 1.07450933e+01 4.03483979e+00-2.15836864e-03 1.18233875e-05    3
-1.18459406e-08 4.00593954e-12 3.83636392e+03 4.20008770e+00                   4
HO2CHO                  C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230825e+01 4.43559488e-03-1.56185338e-06 2.43413972e-10-1.38379570e-14    2
-3.81313380e+04-2.33591553e+01 2.47434345e+00 2.16898555e-02-1.63512196e-05    3
 5.87745825e-09-8.18701426e-13-3.54892793e+04 1.72835404e+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473661e+00 8.42765725e-03-3.84722250e-06 8.63389842e-10-7.73674422e-14    2
-4.73118221e+04 5.12933885e+00 1.85206266e+00 1.27447105e-02-7.44476686e-06    3
 2.19581368e-09-2.62426309e-13-4.66124595e+04 1.56434956e+01                   4
OCHO                    C   1O   2H   1     G    200.00   3500.00  700.00      1
 2.58373953e+00 8.99565940e-03-4.55939787e-06 1.11902584e-09-1.07899898e-13    2
-1.67164582e+04 1.34890938e+01 4.25809175e+00-5.72067562e-04 1.59428742e-05    3
-1.84069475e-08 6.86566202e-12-1.69508675e+04 6.00851172e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959141e+00 1.57445261e-02-5.96197393e-06 1.06867182e-09-7.61012340e-14    2
-1.25948053e+04-1.43089412e+00-2.41778724e-01 2.53475709e-02-1.39645112e-05    3
 4.03257452e-09-4.87754387e-13-1.10391121e+04 2.19572625e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791360e+00 1.11042800e-02-3.71281686e-06 5.47665571e-10-2.89412604e-14    2
 1.17176215e+04-4.91382513e+00 6.75421801e-01 2.11542617e-02-1.20878017e-05    3
 3.64951180e-09-4.59753237e-13 1.33457186e+04 1.95628439e+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   3500.00 1450.00      1
 1.00876750e+01 1.40221806e-02-4.79128015e-06 7.15474133e-10-3.78163629e-14    2
-2.40669299e+04-2.56733582e+01-5.77204918e-01 4.34425389e-02-3.52261336e-05    3
 1.47085102e-08-2.45040879e-12-2.09741147e+04 2.97412031e+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   3500.00 1480.00      1
 9.29919683e+00 1.29334624e-02-4.54028592e-06 7.01327861e-10-3.92078228e-14    2
-7.64002445e+03-2.14311736e+01 2.00183268e-01 3.75253910e-02-2.94645378e-05    3
 1.19284684e-08-1.93568426e-12-4.94671644e+03 2.60335034e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402718e+00 9.50595350e-03-3.15129261e-06 4.53052074e-10-2.23949159e-14    2
 3.97229102e+03-3.77420905e+00-6.02932450e-02 2.08133970e-02-1.34307867e-05    3
 4.60638301e-09-6.51687481e-13 5.51151676e+03 2.10642172e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728376e+00 7.47581588e-03-2.58984227e-06 4.05265795e-10-2.35022721e-14    2
 3.38403785e+04 1.51958751e+00 1.23421214e+00 1.56222204e-02-1.10171572e-05    3
 4.27989337e-09-6.91541509e-13 3.46967692e+04 1.68637048e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267454e+00 5.47212830e-03-2.03181542e-06 3.75019116e-10-2.77049062e-14    2
 2.58626597e+04-2.43835921e+00 7.70536907e-01 2.37107998e-02-3.66622044e-05    3
 2.95989761e-08-9.27579255e-12 2.64317975e+04 1.40907683e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788257e+00 4.21328989e-03-1.58936946e-06 2.68739191e-10-1.73346359e-14    2
 6.72874491e+04 5.32512367e+00 4.60873599e+00 1.42766785e-03 8.54158643e-07    3
-6.83903344e-10 1.21940589e-13 6.68801772e+04-1.05894068e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490827e+00 1.39762977e-02-4.67366748e-06 6.82063684e-10-3.47025038e-14    2
-3.18909574e+04-1.38313071e+01-4.22291411e-01 3.35894614e-02-2.32937596e-05    3
 8.53864266e-09-1.27783209e-12-2.94428423e+04 2.70882146e+01                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957255e+00 2.35453825e-02-1.23415273e-05 3.08911893e-09-2.98016648e-13    2
-3.10347953e+03 1.69410913e+01 3.27852943e+00 1.44656289e-02 7.11508755e-06    3
-1.54409905e-08 6.31987957e-12-3.32593350e+03 9.84203392e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479680e+00 1.17471700e-02-4.06239751e-06 6.31554725e-10-3.61645074e-14    2
-6.24418450e+03-9.60110092e+00 1.82077785e+00 2.63431399e-02-1.89562444e-05    3
 7.38613379e-09-1.18490244e-12-4.66716293e+03 1.83437446e+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1500.00      1
 6.63757422e+00 1.19924585e-02-4.07718738e-06 6.22004997e-10-3.47508084e-14    2
-9.66525354e+03-7.65007787e+00 1.23305393e+00 2.64045127e-02-1.84892415e-05    3
 7.02736239e-09-1.10231037e-12-8.04389745e+03 2.06149529e+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   3500.00 1440.00      1
 9.66417632e+00 1.29483231e-02-4.44318337e-06 6.83406482e-10-3.84804393e-14    2
 1.86599132e+03-2.38806241e+01 2.23212418e+00 3.35929124e-02-2.59479639e-05    3
 1.06393234e-08-1.76693824e-12 4.00642234e+03 1.46847781e+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   3500.00 1520.00      1
 6.04215804e+00 1.11433647e-02-3.80167462e-06 5.65226940e-10-2.94248186e-14    2
-9.44151524e+03-1.02352918e+01-2.19672856e+00 3.28246452e-02-2.51976751e-05    3
 9.94943769e-09-1.57288053e-12-6.93689371e+03 3.29622805e+01                   4
C2H3O1-2                C   2H   3O   1     G    200.00   3500.00 1800.00      1
 7.60993625e+00 6.11300596e-03-1.59366937e-06 1.28294159e-10 2.98968068e-15    2
 1.61313302e+04-1.70584528e+01 7.34197746e-02 2.28608204e-02-1.55501814e-05    3
 5.29737268e-09-7.14937891e-13 1.88444761e+04 2.37307466e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195371e+00 1.06589270e-02-3.75190329e-06 6.00731628e-10-3.66603824e-14    2
-2.30621355e+04-8.31408577e+00 9.75916637e-01 2.23167871e-02-1.34667868e-05    3
 4.19883662e-09-5.36397187e-13-2.11735621e+04 2.00785613e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 6.07689016e+00 8.12979339e-03-2.81854999e-06 4.38698307e-10-2.55171837e-14    2
-4.06801047e+03-6.15492453e+00 1.47388064e+00 1.83587034e-02-1.13426417e-05    3
 3.59576931e-09-4.63999267e-13-2.41092705e+03 1.87575232e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703792e+00 7.91358604e-03-2.83605891e-06 4.62112655e-10-2.83231297e-14    2
-1.16170812e+03-8.37157286e+00 7.37868281e-01 2.50454357e-02-2.20135026e-05    3
 1.00031294e-08-1.80836357e-12 3.76389339e+02 2.09962837e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523628e+00 6.46841658e-03-2.33588414e-06 3.83408110e-10-2.36897850e-14    2
-8.05944305e+03-4.61154403e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226119e-09-9.59140718e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420513e+00 3.89116779e-03-1.41168608e-06 2.35668533e-10-1.49424971e-14    2
 1.94026782e+04-4.94089647e+00 3.33028661e+00 1.20351629e-02-1.14247949e-05    3
 5.70731267e-09-1.13618105e-12 2.00087543e+04 7.53650387e+00                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483420e-03 1.65900439e-06-8.55133989e-10 9.82287244e-14    2
-2.73756816e+04-4.36816973e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH2OHCHO                C   2H   4O   2     G    300.00   3500.00 1800.00      1
 8.91045186e+00 9.14305837e-03-2.53718677e-06 2.39203912e-10 8.50819938e-16    2
-4.09945450e+04-1.84179622e+01 1.56305396e+00 2.54706093e-02-1.61434792e-05    3
 5.27857147e-09-6.99061342e-13-3.83494818e+04 2.13476880e+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   3500.00 1570.00      1
 9.97760259e+00 4.26981223e-03-1.12729433e-06 7.37809055e-11 5.98360578e-15    2
-2.96900177e+04-2.75230973e+01 7.08345765e-01 2.78857532e-02-2.36902952e-05    3
 9.65467301e-09-1.51963616e-12-2.67794711e+04 2.13768445e+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319128e-02-1.90892866e-05    3
 5.92848299e-09-7.42884555e-13-1.63833552e+04 6.70139035e+00                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 5.02910657e+00-2.87377519e-02 6.15808970e-05-2.98073518e-08 4.29774802e-12    2
-4.07046731e+04 1.82412181e+01 2.12034974e-07-1.31715123e-09 2.87530013e-12    3
 2.88411189e-08-1.66481344e-11-4.00005982e+04 4.07099930e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849390e-09-3.11411020e-13    2
-2.07588781e+04 1.60124236e+01 4.66126893e+00 9.68655552e-03 1.14715528e-05    3
-1.83003965e-08 7.03409940e-12-2.10634335e+04 6.60518516e+00                   4
C3H8                    C   3H   8          G    300.00   3500.00 1690.00      1
 8.33847007e+00 1.79340922e-02-5.80534981e-06 7.91037708e-10-3.43401227e-14    2
-1.70816233e+04-2.27461799e+01-1.38651266e+00 4.09518028e-02-2.62352705e-05    3
 8.85017800e-09-1.22652064e-12-1.37945792e+04 2.92742161e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1800.00      1
 6.05951251e+00 1.82035621e-02-6.54041321e-06 1.09272144e-09-7.13189353e-14    2
 7.29671818e+03-6.80793083e+00-6.08211221e-01 3.30207259e-02-1.88880497e-05    3
 5.66592015e-09-7.06485424e-13 9.69709872e+03 2.92791809e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1590.00      1
 7.21724982e+00 1.65877265e-02-5.58902439e-06 8.31338515e-10-4.40999325e-14    2
 8.50975633e+03-1.26938767e+01-1.37086178e-01 3.50892007e-02-2.30432453e-05    3
 8.14967015e-09-1.19478101e-12 1.08484352e+04 2.61969991e+01                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755201e+00 1.65820017e-02-6.59972302e-06 1.29512916e-09-1.03784375e-13    2
-3.79456071e+02-1.05616187e+01-8.55987188e-02 3.08112255e-02-1.84574096e-05    3
 5.68686491e-09-7.13747674e-13 1.92567819e+03 2.40935687e+01                   4
C3H5-A                  C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877792e+00 1.04611885e-02-3.15379708e-06 3.85306884e-10-1.26413689e-14    2
 1.71766363e+04-2.28181758e+01-3.57888096e-01 3.27028536e-02-2.40053580e-05    3
 9.07345729e-09-1.37016487e-12 2.00235695e+04 2.42845603e+01                   4
C3H5-S                  C   3H   5          G    300.00   3500.00 1800.00      1
 6.52599516e+00 1.37686655e-02-5.50691342e-06 1.07278366e-09-8.39560017e-14    2
 2.86430050e+04-9.99635700e+00 1.54227621e+00 2.48435965e-02-1.47360226e-05    3
 4.49097224e-09-5.58704416e-13 3.04371438e+04 1.69765696e+01                   4
C3H5-T                  C   3H   5          G    300.00   3500.00  770.00      1
 1.49331935e+00 2.33788729e-02-1.18550710e-05 2.86552470e-09-2.68203790e-13    2
 2.87117775e+04 1.76892214e+01 2.52238869e+00 1.80330581e-02-1.44114618e-06    3
-6.15086046e-09 2.65919399e-12 2.85533009e+04 1.29935191e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079978e+00 1.37589661e-02-5.15319199e-06 9.32421983e-10-6.74695911e-14    2
 7.77376170e+03-2.10036658e+01 9.27196847e-01 3.40908988e-02-2.40959865e-05    3
 8.77622923e-09-1.28545208e-12 1.04088818e+04 2.23747992e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1550.00      1
 9.00938222e+00 1.57632590e-02-5.29374355e-06 7.64253417e-10-3.74126438e-14    2
-1.56669515e+04-2.44960178e+01-1.88321638e+00 4.38731909e-02-3.24969034e-05    3
 1.24645372e-08-1.92455519e-12-1.22902459e+04 3.28282089e+01                   4
CH3CHCHO                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 6.70347362e+00 1.89922318e-02-9.18109977e-06 2.14445657e-09-1.96154637e-13    2
-6.21094363e+03-1.05801331e+01 2.92067498e-01 3.32398010e-02-2.10540741e-05    3
 6.54185446e-09-8.06904344e-13-3.90283743e+03 2.41197343e+01                   4
AC4H7OOH                C   4H   8O   2     G    300.00   3500.00 1660.00      1
 1.22738272e+01 2.55483383e-02-9.81265077e-06 1.82078670e-09-1.35039880e-13    2
-1.24525960e+04-3.36837474e+01 1.60151447e+00 5.12647544e-02-3.30503762e-05    3
 1.11532065e-08-1.54052480e-12-8.90938817e+03 2.32129081e+01                   4
CH3CHCO                 C   3H   4O   1     G    300.00   3500.00 1280.00      1
 6.99681463e+00 1.49445085e-02-6.71568578e-06 1.45955079e-09-1.25293200e-13    2
-1.29366480e+04-1.07908059e+01 1.50068777e+00 3.21199049e-02-2.68431035e-05    3
 1.19425808e-08-2.17276001e-12-1.15296395e+04 1.70816035e+01                   4
AC3H5OOH                C   3H   6O   2     G    298.00   3500.00 1800.00      1
 1.36957657e+01 1.27112963e-02-4.21186263e-06 6.49030109e-10-3.94931202e-14    2
-1.11479407e+04-4.31791016e+01 4.22354618e+00 3.37606729e-02-2.17530098e-05    3
 7.14575129e-09-9.41815506e-13-7.73794171e+03 8.08652616e+00                   4
C3H6OH1-2               C   3H   7O   1     G    300.00   3500.00 1800.00      1
 8.46016352e+00 1.89669003e-02-7.38013554e-06 1.39189577e-09-1.05413394e-13    2
-1.21581707e+04-1.51603324e+01 4.08605477e-01 3.68592515e-02-2.22904282e-05    3
 6.91422639e-09-8.72403758e-13-9.25960980e+03 2.84163793e+01                   4
C3H6OH2-1               C   3H   7O   1     G    300.00   3500.00 1590.00      1
 8.99548234e+00 1.75103792e-02-6.94615357e-06 1.37004323e-09-1.07539337e-13    2
-1.65436320e+04-1.93287236e+01 1.31207693e+00 3.68397010e-02-2.51813628e-05    3
 9.01583327e-09-1.30970758e-12-1.41003090e+04 2.13023225e+01                   4
HOC3H6O2                C   3H   7O   3     G    300.00   3500.00 1480.00      1
 1.24409055e+01 2.15172909e-02-8.97737594e-06 1.82414691e-09-1.48047122e-13    2
-3.10315628e+04-3.23089026e+01 2.93449048e+00 4.72103044e-02-3.50175923e-05    3
 1.35539741e-08-2.12943685e-12-2.82176640e+04 1.72809693e+01                   4
SC3H5OH                 C   3H   6O   1     G    300.00   3500.00 1260.00      1
 7.83167544e+00 1.85990426e-02-7.98421836e-06 1.67672190e-09-1.40411942e-13    2
-2.22362405e+04-1.56369776e+01-5.71229678e-02 4.36428470e-02-3.77982713e-05    3
 1.74513531e-08-3.27029908e-12-2.02482633e+04 2.42451084e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00 1630.00      1
 9.39463114e+00 1.51343106e-02-4.86246276e-06 6.64177249e-10-2.94552530e-14    2
-2.20582199e+04-2.45922026e+01 4.73537667e-01 3.70265645e-02-2.50087087e-05    3
 8.90395064e-09-1.29322418e-12-1.91499434e+04 2.28055845e+01                   4
CH2CCH2OH               C   3H   5O   1     G    300.00   3500.00 1800.00      1
 7.15397365e+00 1.62590933e-02-7.06959971e-06 1.52062107e-09-1.30983749e-13    2
 1.01359982e+04-8.36739478e+00 2.39300609e+00 2.68390212e-02-1.58862063e-05    3
 4.78603091e-09-5.84512894e-13 1.18499465e+04 1.73999548e+01                   4
C3H4-P                  C   3H   4          G    300.00   3500.00 1570.00      1
 6.45797858e+00 1.06371316e-02-3.61161722e-06 5.39412691e-10-2.85851275e-14    2
 1.94136786e+04-1.10770989e+01 1.72714322e+00 2.26902153e-02-1.51273023e-05    3
 5.42930020e-09-8.07229635e-13 2.08991609e+04 1.38804115e+01                   4
C3H4-A                  C   3H   4          G    300.00   3500.00 1420.00      1
 6.37608366e+00 1.10282079e-02-3.89476312e-06 6.16686076e-10-3.59564768e-14    2
 2.00917847e+04-1.13283006e+01 5.08248696e-01 2.75573205e-02-2.13550933e-05    3
 8.81402419e-09-1.47914981e-12 2.17582498e+04 1.90382079e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057762e+00 1.05635747e-02-4.84060952e-06 1.09040068e-09-9.80036130e-14    2
 4.00565408e+04-5.04125059e+00 1.75584147e+00 2.95861278e-02-3.88094543e-05    3
 2.80498013e-08-8.12163476e-12 4.07276565e+04 1.35345464e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00 1260.00      1
 6.42043189e+00 6.05128866e-03-2.30888141e-06 4.10631875e-10-2.84293474e-14    2
 6.08598164e+04-8.32404334e+00 2.15397882e+00 1.95955841e-02-1.84330427e-05    3
 8.94193413e-09-1.72114805e-12 6.19349626e+04 1.32451538e+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1710.00      1
 9.33264604e+00 1.46861072e-02-4.56011955e-06 5.69518135e-10-1.90908109e-14    2
-2.69164882e+04-2.52385565e+01-9.86882752e-02 3.67477080e-02-2.39124009e-05    3
 8.11426720e-09-1.12212430e-12-2.36909719e+04 2.53220280e+01                   4
CH2CH2CHO               C   3H   5O   1     G    300.00   3500.00  700.00      1
 1.38640400e+00 2.84363938e-02-1.56688640e-05 4.07196321e-09-4.03232083e-13    2
 6.14151634e+02 2.19844218e+01 2.41071832e+00 2.25831692e-02-3.12623980e-06    3
-7.87339320e-09 3.86296664e-12 4.70747631e+02 1.74080446e+01                   4
RALD3                   C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180078e-02-2.61696720e-05 6.65382129e-09-6.35305357e-13    2
-2.14966001e+03 5.90959840e+01 7.04072886e+00-2.01204450e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381685e+00                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597839e+00 1.12038372e-02-3.67974365e-06 5.08180252e-10-2.25803375e-14    2
-1.23719484e+04-2.08137560e+01 8.18908043e-01 3.22215131e-02-2.33838148e-05    3
 8.71820989e-09-1.30539747e-12-9.68168587e+03 2.36968522e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00 1790.00      1
 9.79507855e+00 1.35932465e-02-4.01642284e-06 4.43034305e-10-7.94380246e-15    2
-3.07542949e+04-2.70699391e+01-7.54581368e-03 3.54985524e-02-2.23728244e-05    3
 7.27968292e-09-9.62782995e-13-2.72449554e+04 2.59292980e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1590.00      1
 8.40473847e+00 1.29432044e-02-4.25667366e-06 6.02254911e-10-2.86748418e-14    2
-7.89528923e+03-1.63899805e+01 1.00367440e+00 3.15622335e-02-2.18217955e-05    3
 7.96708586e-09-1.18666713e-12-5.54175085e+03 2.27480006e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14851999e-06-5.94424210e-11 5.32964638e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
PC4H9                   C   4H   9          G    300.00   3500.00  950.00      1
 3.94763006e+00 3.16286394e-02-1.12984867e-05 1.11637450e-09 5.54031605e-14    2
 6.05554723e+03 7.76350061e+00-2.76188385e-01 4.94131381e-02-3.93792741e-05    3
 2.08221903e-08-5.13033783e-12 6.85807273e+03 2.79243295e+01                   4
SC4H9                   C   4H   9          G    300.00   3500.00  850.00      1
 3.40122928e+00 3.20901863e-02-1.12255470e-05 9.71712110e-10 8.30726274e-14    2
 4.66283101e+03 1.05291639e+01 2.36336421e-01 4.69837998e-02-3.75083943e-05    3
 2.15857099e-08-5.97986791e-12 5.20086280e+03 2.52835874e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955795e+00 3.23747266e-02-1.18655436e-05 1.37455177e-09 1.57073481e-14    2
-1.97025810e+04-6.34483426e+00-1.85965329e+00 5.58007941e-02-3.97537191e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H9                   C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221490e-06 8.09648920e-10 4.02033223e-14    2
 3.37759297e+03-1.61084037e+01-1.15582377e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
TC4H9                   C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871689e+00 2.55264450e-02-8.65284049e-06 8.24419700e-10 3.80550657e-14    2
 8.35470579e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397361e-05    3
 1.42467509e-08-2.35878980e-12 3.41363196e+03 3.01901373e+01                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385767e+03-1.72949366e+01 7.17301599e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035733e-13-3.72372397e+03 2.01415164e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177117e+00 3.67769037e-02-1.77031337e-05 3.74786266e-09-2.92191284e-13    2
 1.31214242e+04 2.00120540e+01 3.86130010e+00 2.14653098e-02 1.51074247e-05    3
-2.75002882e-08 1.08678626e-11 1.27462902e+04 8.04059663e+00                   4
IC4H7O                  C   4H   7O   1     G    300.00   3500.00 1800.00      1
 1.18822163e+01 1.89918532e-02-7.42296498e-06 1.41442848e-09-1.08683660e-13    2
 1.15971319e+03-3.56333819e+01 1.50010972e+00 4.20632012e-02-2.66490883e-05    3
 8.53521488e-09-1.09768177e-12 4.89727156e+03 2.05567447e+01                   4
C4H8-1                  C   4H   8          G    300.00   3500.00 1800.00      1
 1.03330449e+01 1.99470428e-02-7.40538998e-06 1.30472507e-09-9.09598189e-14    2
-5.56551437e+03-3.07722296e+01-6.91489888e-01 4.44460090e-02-2.78211951e-05    3
 8.86613439e-09-1.14115556e-12-1.59668184e+03 2.88948525e+01                   4
C4H8-2                  C   4H   8          G    300.00   3500.00 1800.00      1
 5.15907399e+00 2.89997694e-02-1.32974598e-05 2.96139017e-09-2.60424474e-13    2
-4.76704683e+03-3.39008062e+00 5.60608454e-01 3.92185817e-02-2.18131368e-05    3
 6.11534459e-09-6.98473698e-13-3.11159924e+03 2.14977742e+01                   4
C4H71-3                 C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017754e+00 1.98466503e-02-6.37614061e-06 5.28652768e-10 3.81103734e-14    2
 1.19533850e+04-1.83767119e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
C4H71-4                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075605e-06 3.82147970e-10 5.73994809e-14    2
 1.98988324e+04-1.80212793e+01-3.29329052e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
C4H71-O                 C   4H   7O   1     G    300.00   3500.00 1600.00      1
 1.37371777e+01 1.70982846e-02-6.55972544e-06 1.21466090e-09-8.98269615e-14    2
-3.28789072e+01-4.64105970e+01-1.48200925e+00 5.51462520e-02-4.22296948e-05    3
 1.60771481e-08-2.41209059e-12 4.83726091e+03 3.41662556e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872521e+00 1.50139591e-02-5.06688177e-06 7.84148097e-10-4.70262839e-14    2
 8.60829987e+03-2.47389586e+01 4.65225109e-01 3.46661815e-02-2.14437338e-05    3
 6.84964885e-09-8.89456944e-13 1.17919599e+04 2.31239087e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794386e-03 4.88814514e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742308e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777119e+00 1.26498258e-02-4.62248950e-06 7.81217082e-10-5.07629107e-14    2
 3.13366016e+04-1.49692661e+01 7.13119716e-01 3.41836288e-02-2.96617954e-05    3
 1.37214268e-08-2.55855550e-12 3.31283217e+04 2.03030643e+01                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590364e-03 1.80568200e-06-9.30237204e-10 1.18077198e-13    2
 6.01811751e+04-4.25791500e+01 2.34662666e+00 2.83894138e-02-2.35278181e-05    3
 9.69177543e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00  720.00      1
 7.13414735e+00 1.00526308e-02-4.84819206e-06 1.14884604e-09-1.07722834e-13    2
 5.27577824e+04-1.36443516e+01-4.34754087e-01 5.21020832e-02-9.24512179e-05    3
 8.22627589e-08-2.82722759e-11 5.38477042e+04 2.03848077e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055544e+01 1.99961045e-02-7.07935460e-06 1.10673028e-09-6.24178899e-14    2
 4.11452290e+03-4.24445091e+01-6.99882110e+00 7.24907868e-02-6.29247613e-05    3
 2.75111779e-08-4.74405754e-12 9.33275680e+03 5.31863191e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152220e+01 1.47750067e-02-3.90939181e-06 2.82308156e-10 1.62511622e-14    2
 1.91167581e+04-5.54965184e+01-3.67012639e+00 6.11476948e-02-4.84985149e-05    3
 1.93374890e-08-3.03746371e-12 2.47593868e+04 3.97971310e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331261e+01 1.77269649e-02-6.33615682e-06 1.00236865e-09-5.75481750e-14    2
 3.49856300e+04-3.80075865e+01-6.76261385e+00 6.95132669e-02-6.22206553e-05    3
 2.78054854e-08-4.87825263e-12 3.99884457e+04 5.47375207e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786764e+01 1.28174257e-02-3.11961936e-06 1.29368393e-10 2.76958521e-14    2
 9.43770579e+03-5.26289052e+01-4.05866643e+00 5.60992486e-02-4.29495178e-05    3
 1.64197154e-08-2.47082363e-12 1.51874796e+04 4.10783319e+01                   4
C5H5                    H   5C   5          G    200.00   3500.00 1290.00      1
 6.86396822e+00 2.31427769e-02-1.13257692e-05 2.70799252e-09-2.56251711e-13    2
 2.77724452e+04-1.52693149e+01-3.43772279e+00 5.50860048e-02-4.84690575e-05    3
 2.19034903e-08-3.97630943e-12 3.04302815e+04 3.70536347e+01                   4
C5H5CH3                 C   6H   8          G    300.00   3500.00 1470.00      1
 1.21408016e+01 2.34281374e-02-7.98702759e-06 1.18908391e-09-6.20202054e-14    2
 7.23040214e+03-4.21606537e+01-5.49894699e+00 7.14274534e-02-5.69659215e-05    3
 2.34017342e-08-3.83968182e-12 1.24164882e+04 4.97368686e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248658e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987877e+01                   4
C5H5OH                  C   5H   6O   1     G    200.00   3500.00 1450.00      1
 1.34279261e+01 1.64213103e-02-5.21419394e-06 6.78762290e-10-2.54882777e-14    2
-1.08112826e+04-4.76154890e+01-3.54477524e+00 6.32425554e-02-5.36499648e-05    3
 2.29480822e-08-3.86502620e-12-5.88919918e+03 4.05744212e+01                   4
C5H5O                   H   5C   5O   1     G    200.00   3500.00 1380.00      1
 7.52425952e+00 2.65795845e-02-1.33939818e-05 3.28296341e-09-3.17054855e-13    2
 4.64512525e+02-1.52910629e+01-2.58346517e+00 5.58773372e-02-4.52393652e-05    3
 1.86672066e-08-3.10405543e-12 3.25424454e+03 3.67283973e+01                   4
C5H4OH                  H   5C   5O   1     G    200.00   3500.00 1290.00      1
 8.68429815e+00 2.48368249e-02-1.26118784e-05 3.11347632e-09-3.02421966e-13    2
 3.90640044e+03-2.17291570e+01-3.25514699e+00 6.18583602e-02-5.56601753e-05    3
 2.53606582e-08-4.61389132e-12 6.98677728e+03 3.89120509e+01                   4
C5H4O                   C   5H   4O   1     G    200.00   3500.00 1550.00      1
 1.18776174e+01 1.30371391e-02-3.92696670e-06 4.38039798e-10-7.33842917e-15    2
 1.13417720e+03-3.96157060e+01-1.34835256e+00 4.71686744e-02-3.69574847e-05    3
 1.46447142e-08-2.29873753e-12 5.23422788e+03 2.99883001e+01                   4
NC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1650.00      1
 9.25591855e+00 2.27563801e-02-9.54934453e-06 1.92559465e-09-1.53946670e-13    2
-9.34005086e+03-1.86388081e+01 1.92964396e+00 4.05170458e-02-2.56954042e-05    3
 8.44925513e-09-1.14238008e-12-6.92238025e+03 2.03750491e+01                   4
IC3H7O2                 C   3H   7O   2     G    300.00   3500.00 1260.00      1
 7.34738699e+00 2.68252330e-02-1.24179691e-05 2.76645854e-09-2.42147350e-13    2
-1.06484855e+04-8.92587195e+00 1.07341266e+00 4.67426118e-02-3.61291344e-05    3
 1.53120486e-08-2.73135173e-12-9.06744395e+03 2.27924165e+01                   4
C3H7OOH                 C   3H   8O   2     G    300.00   3500.00 1530.00      1
 1.13871492e+01 1.97925480e-02-6.62893779e-06 9.67106876e-10-4.94700798e-14    2
-2.73563036e+04-2.91104777e+01-9.73590405e-01 5.21082072e-02-3.83109566e-05    3
 1.47719081e-08-2.30515656e-12-2.35739173e+04 3.57795697e+01                   4
C3-OQOOH                C   3H   6O   3     G    300.00   3500.00 1350.00      1
 1.12132537e+01 2.34709018e-02-1.13098317e-05 2.59008079e-09-2.30885269e-13    2
-3.91289882e+04-2.66260028e+01 8.46220450e-01 5.41880374e-02-4.54399823e-05    3
 1.94444762e-08-3.35206960e-12-3.63298893e+04 2.65001343e+01                   4
CHOCH2CHO               C   3H   4O   2     G    300.00   3500.00 1370.00      1
 1.06304440e+01 1.18394227e-02-4.21486308e-06 6.67473434e-10-3.88516159e-14    2
-4.37970340e+04-2.83088260e+01-8.46550190e-01 4.53488948e-02-4.09040660e-05    3
 1.85211002e-08-3.29681270e-12-4.06523375e+04 3.06741176e+01                   4
CH2OHCH2CHO             C   3H   6O   2     G    300.00   3500.00 1800.00      1
 1.08721654e+01 1.63593216e-02-6.08637842e-06 1.10130849e-09-8.02911325e-14    2
-4.55272952e+04-2.70748520e+01 2.66105929e+00 3.46062241e-02-2.12921305e-05    3
 6.73306853e-09-8.62480026e-13-4.25712970e+04 1.73653673e+01                   4
CH3CO2H                 C   2H   4O   2     G    300.00   3500.00 1800.00      1
 1.06195365e+01 8.83226600e-03-2.54924379e-06 2.13473353e-10 7.27652554e-15    2
-5.71972759e+04-3.23726793e+01-7.52613551e-01 3.41037106e-02-2.36087809e-05    3
 8.01330193e-09-1.07603300e-12-5.31033019e+04 2.91757692e+01                   4
HCO3                    C   1H   1O   3     G    300.00   3500.00 1490.00      1
 7.67843584e+00 4.62692543e-03-1.54275270e-06 2.12409842e-10-8.98166116e-15    2
-1.61147276e+04-1.27152259e+01 2.31459990e+00 1.90264850e-02-1.60389536e-05    3
 6.69840577e-09-1.09723601e-12-1.45163044e+04 1.53011516e+01                   4
HCO3H                   C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230668e+01 4.43563253e-03-1.56188514e-06 2.43424395e-10-1.38391380e-14    2
-3.81313332e+04-2.33590722e+01 2.47434199e+00 2.16898607e-02-1.63512235e-05    3
 5.87745807e-09-8.18701091e-13-3.54892796e+04 1.72835470e+01                   4
CH2OHCOCH3              C   3H   6O   2     G    300.00   3500.00 1460.00      1
 1.16062110e+01 1.59761333e-02-5.42430575e-06 8.11522092e-10-4.31363774e-14    2
-4.81919050e+04-3.20429615e+01 9.15361352e-01 4.52661324e-02-3.55167705e-05    3
 1.45523736e-08-2.39602191e-12-4.50701769e+04 2.35800153e+01                   4
NC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1800.00      1
 1.29748618e+01 1.76433870e-02-7.16935406e-06 1.42696153e-09-1.14477043e-13    2
-5.86411825e+03-3.67690498e+01 1.55643299e+00 4.30176732e-02-2.83145926e-05    3
 9.25853134e-09-1.20219507e-12-1.75348388e+03 2.50298688e+01                   4
IC3-QOOH                C   3H   7O   2     G    300.00   3500.00 1270.00      1
 1.04498043e+01 2.29490980e-02-1.05757759e-05 2.34172678e-09-2.03669154e-13    2
-5.22299426e+03-2.40008692e+01-1.71110877e-01 5.64007993e-02-5.00856593e-05    3
 2.30818230e-08-4.28636527e-12-2.52528181e+03 2.97774852e+01                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1260.00      1
 1.11683562e+01 2.95822139e-02-1.42526305e-05 3.27126849e-09-2.92476812e-13    2
-2.00281219e+04-2.06289848e+01 2.57588692e+00 5.68598942e-02-4.67260594e-05    3
 2.04529769e-08-3.70154594e-12-1.78628196e+04 2.28105329e+01                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   3500.00 1220.00      1
 1.23035624e+01 2.79964884e-02-1.33482910e-05 3.03524084e-09-2.69271163e-13    2
-2.25784829e+04-2.78550798e+01 1.73143844e+00 6.26591899e-02-5.59663668e-05    3
 2.63238068e-08-5.04151829e-12-1.99988847e+04 2.52515831e+01                   4
CH2COOH                 C   2H   3O   2     G    300.00   3500.00 1440.00      1
 1.01170850e+01 5.56298782e-03-8.24128628e-07-2.50442742e-11 1.25384218e-14    2
-3.40138321e+04-2.77197730e+01 4.26277933e-01 3.24818963e-02-2.88646583e-05    3
 1.29566824e-08-2.24123357e-12-3.12228797e+04 2.25664553e+01                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1570.00      1
 1.51567879e+01 2.57227734e-02-1.11020451e-05 2.28943518e-09-1.86269530e-13    2
-4.30658407e+04-4.59845002e+01 9.69279338e-01 6.18692920e-02-4.56369355e-05    3
 1.69539322e-08-2.52138051e-12-3.86109630e+04 2.88616666e+01                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   3500.00 1330.00      1
 1.18153445e+01 3.20093755e-02-1.53334982e-05 3.50316407e-09-3.12136547e-13    2
-4.27660549e+04-2.73083214e+01 2.51946601e+00 5.99669047e-02-4.68645461e-05    3
 1.93082006e-08-3.28300808e-12-4.02933512e+04 2.01899074e+01                   4
C4H9OOH                 C   4H  10O   2     G    300.00   3500.00 1780.00      1
 1.73966948e+01 2.30088698e-02-8.34646932e-06 1.39883190e-09-9.01677554e-14    2
-3.38614042e+04-6.23628946e+01 1.12895120e+00 5.95655969e-02-3.91527000e-05    3
 1.29367460e-08-1.71066131e-12-2.80700874e+04 2.54997628e+01                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   3500.00 1580.00      1
 1.69833146e+01 2.73095032e-02-1.19226853e-05 2.48166925e-09-2.03420392e-13    2
-3.51234520e+04-5.58041780e+01 1.44561329e+00 6.66454559e-02-4.92669442e-05    3
 1.82387405e-08-2.69662788e-12-3.02135384e+04 2.62635800e+01                   4
NC5H10-O                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.40073101e+01 3.04405284e-02-1.35854526e-05 2.90305354e-09-2.44985844e-13    2
-2.55455866e+04-5.25239383e+01-3.79263098e+00 6.99959530e-02-4.65483064e-05    3
 1.51115179e-08-1.94060590e-12-1.91376078e+04 4.38130562e+01                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   3500.00 1410.00      1
 1.42172630e+01 3.77707683e-02-1.76257936e-05 3.93443034e-09-3.43954252e-13    2
-4.65061050e+04-3.85369191e+01 2.52749929e+00 7.09332187e-02-5.29049961e-05    3
 2.06149043e-08-3.30148510e-12-4.32095916e+04 2.18759162e+01                   4
NC5H11OOH               C   5H  12O   2     G    300.00   3500.00 1630.00      1
 1.66988185e+01 3.44172712e-02-1.43139761e-05 2.85300849e-09-2.25350876e-13    2
-3.73755763e+04-5.75775302e+01 6.24289379e-02 7.52427671e-02-5.18834508e-05    3
 1.82188468e-08-2.58207455e-12-3.19521133e+04 3.08116402e+01                   4
NC4-QOOH                C   4H   9O   2     G    300.00   3500.00 1760.00      1
 1.83774568e+01 1.83354725e-02-6.23923380e-06 9.66797423e-10-5.61281944e-14    2
-1.29135491e+04-6.55986639e+01 1.19976578e+00 5.73756794e-02-3.95121374e-05    3
 1.35701700e-08-1.84637998e-12-6.86700189e+03 2.69845517e+01                   4
NC4H9-OO                C   4H   9O   2     G    300.00   3500.00 1320.00      1
 8.96630114e+00 3.41074657e-02-1.57641000e-05 3.50715782e-09-3.06662916e-13    2
-1.40847395e+04-1.58347447e+01 9.44281656e-01 5.84166156e-02-4.33881341e-05    3
 1.74586902e-08-2.94899859e-12-1.19669263e+04 2.50940293e+01                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   3500.00 1260.00      1
 9.11667611e+00 3.41757258e-02-1.58797345e-05 3.54686464e-09-3.10976548e-13    2
-1.64591648e+04-1.96564028e+01 4.84069010e-01 6.15808277e-02-4.85048558e-05    3
 2.08088336e-08-3.73597039e-12-1.42837478e+04 2.39860330e+01                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   3500.00 1270.00      1
 1.20890742e+01 3.03954175e-02-1.40883982e-05 3.13822121e-09-2.74437748e-13    2
-1.09705556e+04-3.28537329e+01-4.26302142e-01 6.98139255e-02-6.06456912e-05    3
 2.75777451e-08-5.08536764e-12-7.79165002e+03 3.05171096e+01                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   3500.00 1350.00      1
 1.14809469e+01 3.08095616e-02-1.41939360e-05 3.14755455e-09-2.74422165e-13    2
-7.45268236e+03-2.80879239e+01-1.93281563e-01 6.53998681e-02-5.26276099e-05    3
 2.21271466e-08-3.78916143e-12-4.30064068e+03 3.17369695e+01                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   3500.00 1380.00      1
 8.54295826e+00 3.45220773e-02-1.59311943e-05 3.53852672e-09-3.08950056e-13    2
-1.29532173e+04-1.39825068e+01 7.00555203e-01 5.72536803e-02-4.06394585e-05    3
 1.54748862e-08-2.47133403e-12-1.07887140e+04 2.63784632e+01                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   3500.00 1230.00      1
 1.51474113e+01 3.37812811e-02-1.58996825e-05 3.57608795e-09-3.14486518e-13    2
-2.85698876e+04-4.24732202e+01 1.10123476e+00 7.94599040e-02-7.16053202e-05    3
 3.37688455e-08-6.45122585e-12-2.51145282e+04 2.81992196e+01                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1240.00      1
 1.39939782e+01 3.54845223e-02-1.68915059e-05 3.83671077e-09-3.40131615e-13    2
-2.83614519e+04-3.70531088e+01 1.55094394e+00 7.56233423e-02-6.54465302e-05    3
 2.99415625e-08-5.60320657e-12-2.52755794e+04 2.56539769e+01                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   3500.00 1290.00      1
 1.30518446e+01 3.65484801e-02-1.74274782e-05 3.96741951e-09-3.52552034e-13    2
-2.47096139e+04-3.04334702e+01 1.64511787e+00 7.19181753e-02-5.85550308e-05    3
 2.52219687e-08-4.47165071e-12-2.17666784e+04 2.75020267e+01                   4
C5EN-QOOH               C   5H   9O   2     G    300.00   3500.00 1420.00      1
 1.28791275e+01 3.32930454e-02-1.55378924e-05 3.46674396e-09-3.02869803e-13    2
 3.23011716e+03-3.38507184e+01 1.34404411e+00 6.57862381e-02-4.98616876e-05    3
 1.95812018e-08-3.13992224e-12 6.50608085e+03 2.58442475e+01                   4
C5EN-OO                 C   5H   9O   2     G    300.00   3500.00 1280.00      1
 1.00840321e+01 3.69913036e-02-1.74216180e-05 3.93130749e-09-3.47257402e-13    2
-8.98415155e+02-1.96513637e+01 4.09897282e-01 6.72229749e-02-5.28493577e-05    3
 2.23832553e-08-3.95115346e-12 1.57816336e+03 2.94089022e+01                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   3500.00 1160.00      1
 1.36699765e+01 4.21231934e-02-2.15503712e-05 5.21806335e-09-4.87293013e-13    2
-1.42354804e+04-3.35883365e+01 5.24578569e-01 8.74521518e-02-8.01654036e-05    3
 3.89048636e-08-7.74737927e-12-1.11857480e+04 3.17816498e+01                   4
NC5H12OO                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.06544848e+01 4.16170555e-02-1.93382868e-05 4.32113942e-09-3.79088223e-13    2
-1.98652039e+04-2.50234586e+01 3.19664881e-01 7.34165014e-02-5.60299551e-05    3
 2.31373796e-08-3.99759595e-12-1.71781508e+04 2.75475609e+01                   4
NC5-QOOH                C   5H  11O   2     G    300.00   3500.00 1300.00      1
 1.36538194e+01 3.77860020e-02-1.75151081e-05 3.90394425e-09-3.41708560e-13    2
-1.43879859e+04-3.94678820e+01-5.74283056e-01 8.15647789e-02-6.80290814e-05    3
 2.98085460e-08-5.32336273e-12-1.06886793e+04 3.29074336e+01                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   3500.00 1270.00      1
 1.54638476e+01 4.30531975e-02-2.04284728e-05 4.63174721e-09-4.10271992e-13    2
-3.17413365e+04-4.31406916e+01 1.43265567e+00 8.72459280e-02-7.26246112e-05    3
 3.20312949e-08-5.80388375e-12-2.81774138e+04 2.79053907e+01                   4
C4H6O2                  C   4H   6O   2     G    300.00   3500.00 1800.00      1
 7.01919581e+00 2.89919962e-02-1.39811163e-05 3.22750474e-09-2.90888809e-13    2
-4.36055710e+04-7.47846941e+00 9.15158242e-01 4.25565241e-02-2.52848896e-05    3
 7.41408744e-09-8.72358628e-13-4.14081175e+04 2.55578553e+01                   4
C4H8O                   C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.12815996e+01 2.48463701e-02-1.13234700e-05 2.47069946e-09-2.12413507e-13    2
-2.03756688e+04-3.84267373e+01-2.94845122e+00 5.64687053e-02-3.76754160e-05    3
 1.22306795e-08-1.56796629e-12-1.52528505e+04 3.85892666e+01                   4
C5H8O                   C   5H   8O   1     G    300.00   3500.00 1330.00      1
 6.70800689e+00 3.65243774e-02-1.77765821e-05 4.15639147e-09-3.79163308e-13    2
-5.52771783e+03-9.67918423e+00-5.12640161e+00 7.21165835e-02-5.79181679e-05    3
 2.42774871e-08-4.16132414e-12-2.37976516e+03 5.07899200e+01                   4
RNC3OHOOX               C   3H   7O   3     G    300.00   3500.00 1800.00      1
 3.74667463e+01 1.57251521e-02-1.09732359e-05 3.61008695e-09-4.15087643e-13    2
-5.05275840e+04-1.70384641e+02-4.06427158e+00 1.08016303e-01-8.78825284e-05    3
 3.20950101e-08-4.37132697e-12-3.55764175e+04 5.43898920e+01                   4
QNC3OHOOX               C   3H   7O   3     G    300.00   3500.00 1800.00      1
 3.65507236e+01 1.64042711e-02-1.14786982e-05 3.72939657e-09-4.24702220e-13    2
-4.45414828e+04-1.61156347e+02-1.59743882e+00 1.01177965e-01-8.21234434e-05    3
 2.98941170e-08-4.05869117e-12-3.08081443e+04 4.53094659e+01                   4
ZNC3OHOOX               C   3H   7O   5     G    300.00   3500.00 1140.00      1
 2.54947978e+01 2.87030586e-02-3.65256136e-06-1.12208479e-09 2.39300453e-13    2
-5.46882917e+04-8.79716227e+01-1.83124940e+00 1.24583926e-01-1.29811597e-04    3
 7.26551292e-08-1.59399131e-11-4.84579529e+04 4.74412435e+01                   4
KEHYNC3OH               C   3H   6O   4     G    300.00   3500.00  990.00      1
 2.03864541e+01 2.59482570e-02 2.17638828e-06-3.94711666e-09 6.27440484e-13    2
-7.09480080e+04-6.09332091e+01-1.73111577e+00 1.15312176e-01-1.33223488e-04    3
 8.72312515e-08-2.23973999e-11-6.65687291e+04 4.55489913e+01                   4
C3OHCYETH               C   3H   6O   2     G    200.00   3500.00 1670.00      1
 1.35374623e+01 1.18925361e-02-2.94432280e-06 1.64020760e-10 1.84651199e-14    2
-3.51827731e+04-4.61976551e+01-8.63499032e-01 4.63858566e-02-3.39263472e-05    3
 1.25320944e-08-1.83304291e-12-3.03728520e+04 3.06638119e+01                   4
RBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1670.00      1
 1.45390319e+01 2.69797332e-02-1.09312485e-05 2.12602294e-09-1.64284673e-13    2
-3.56893368e+04-4.22613629e+01 3.26237571e+00 5.39896881e-02-3.51916871e-05    3
 1.18108288e-08-1.61410590e-12-3.19229337e+04 1.79249204e+01                   4
QBU1OOX                 C   4H   9O   3     G    300.00   3500.00 1270.00      1
 9.44680464e+00 1.40890825e-02-6.70668583e-06 1.51288685e-09-1.32818575e-13    2
 1.91332917e+04-2.81812928e+01-5.88861872e+00 6.23896285e-02-6.37545748e-05    3
 3.14592853e-08-6.02777890e-12 2.30284892e+04 4.94686856e+01                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   3500.00 1410.00      1
 1.71509971e+01 3.21642995e-02-1.45265250e-05 3.16055984e-09-2.71089893e-13    2
-4.87167967e+04-4.94521678e+01 4.90929016e+00 6.68925461e-02-5.14714682e-05    3
 2.06286181e-08-3.36826334e-12-4.52646353e+04 1.38131161e+01                   4
KEHYBU1                 C   4H   8O   4     G    300.00   3500.00 1200.00      1
 1.50812003e+01 2.99746636e-02-1.37944087e-05 3.03171374e-09-2.60935207e-13    2
-6.34178095e+04-4.27051070e+01-4.53521778e+00 9.53627237e-02-9.55294839e-05    3
 4.84400889e-08-9.72101336e-12-5.87098692e+04 5.55092666e+01                   4
C4OHCYETH               C   4H   8O   2     G    300.00   3500.00 1740.00      1
 1.55057879e+01 1.98739172e-02-6.85214253e-06 1.07267979e-09-6.29459284e-14    2
-5.34275304e+04-5.89096440e+01-4.24192760e+00 6.52709644e-02-4.59875281e-05    3
 1.60670804e-08-2.21731383e-12-4.65553254e+04 4.72996339e+01                   4
RPENT1OOX               C   5H  11O   3     G    300.00   3500.00 1690.00      1
 2.06735965e+01 3.07535003e-02-1.19967966e-05 2.22747934e-09-1.63728823e-13    2
-5.79272409e+04-7.43003206e+01 2.17872347e+00 7.45283477e-02-5.08502115e-05    3
 1.75542702e-08-2.43100558e-12-5.16759738e+04 2.46315384e+01                   4
QPENT1OOX               C   5H  11O   3     G    300.00   3500.00 1590.00      1
 1.99691781e+01 3.07316205e-02-1.29590658e-05 2.61520663e-09-2.08804310e-13    2
-3.62027680e+04-6.96874635e+01 1.91284982e+00 7.61563458e-02-5.58125803e-05    3
 2.05831372e-08-3.03395063e-12-3.04608556e+04 2.57972168e+01                   4
ZPENT1OOX               C   5H  11O   5     G    300.00   3500.00 1380.00      1
 2.07046201e+01 3.73731215e-02-1.71331760e-05 3.77821832e-09-3.27723702e-13    2
-5.43479695e+04-6.52594396e+01 3.53770719e+00 8.71322894e-02-7.12192280e-05    3
 2.99067459e-08-5.06115261e-12-4.96099015e+04 2.30901712e+01                   4
KEHYP1OH                C   5H  10O   4     G    300.00   3500.00 1560.00      1
 1.98034553e+01 3.06181827e-02-1.26872575e-05 2.52829428e-09-2.00061891e-13    2
-6.77003656e+04-6.61563411e+01 2.43438019e+00 7.51542727e-02-5.55104210e-05    3
 2.08287915e-08-3.13283388e-12-6.22812142e+04 2.53631875e+01                   4
C5OHCYETH               C   5H  10O   2     G    300.00   3500.00 1760.00      1
 1.88847135e+01 2.52072188e-02-8.75962855e-06 1.38787301e-09-8.30558164e-14    2
-5.99419469e+04-8.09815573e+01-5.15784754e+00 7.98494029e-02-5.53296718e-05    3
 1.90280409e-08-2.58876148e-12-5.14789654e+04 4.86014934e+01                   4
RC6OHOOX                C   6H  13O   3     G    300.00   3500.00 1800.00      1
 3.74667463e+01 1.57251521e-02-1.09732359e-05 3.61008695e-09-4.15087643e-13    2
-5.05275840e+04-1.70384641e+02-4.06427158e+00 1.08016303e-01-8.78825284e-05    3
 3.20950101e-08-4.37132697e-12-3.55764175e+04 5.43898920e+01                   4
QC6OHOOX                C   6H  13O   3     G    300.00   3500.00 1800.00      1
 3.65507236e+01 1.64042711e-02-1.14786982e-05 3.72939657e-09-4.24702220e-13    2
-4.45414828e+04-1.61156347e+02-1.59743882e+00 1.01177965e-01-8.21234434e-05    3
 2.98941170e-08-4.05869117e-12-3.08081443e+04 4.53094659e+01                   4
ZC6OHOOX                C   6H  13O   5     G    300.00   3500.00 1140.00      1
 2.54947978e+01 2.87030586e-02-3.65256136e-06-1.12208479e-09 2.39300453e-13    2
-5.46882917e+04-8.79716227e+01-1.83124940e+00 1.24583926e-01-1.29811597e-04    3
 7.26551292e-08-1.59399131e-11-4.84579529e+04 4.74412435e+01                   4
KEHYC6OH                C   6H  12O   4     G    300.00   3500.00  990.00      1
 2.03864541e+01 2.59482570e-02 2.17638828e-06-3.94711666e-09 6.27440484e-13    2
-7.09480080e+04-6.09332091e+01-1.73111577e+00 1.15312176e-01-1.33223488e-04    3
 8.72312515e-08-2.23974000e-11-6.65687291e+04 4.55489913e+01                   4
C6OHCYETH               C   6H  12O   2     G    300.00   3500.00 1760.00      1
 1.88847135e+01 2.52072188e-02-8.75962855e-06 1.38787301e-09-8.30558164e-14    2
-5.99419469e+04-8.09815573e+01-5.15784754e+00 7.98494029e-02-5.53296718e-05    3
 1.90280409e-08-2.58876148e-12-5.14789654e+04 4.86014934e+01                   4
RALD3OO                 C   3H   5O   3     G    300.00   3500.00 1800.00      1
 1.58771657e+01 1.28699615e-02-5.29703385e-06 1.04001953e-09-8.12487153e-14    2
-2.38887629e+04-5.44666587e+01 3.38301196e+00 4.06347476e-02-2.84343556e-05    3
 9.60939795e-09-1.27144016e-12-1.93908676e+04 1.31543077e+01                   4
QALD3OO                 C   3H   5O   3     G    300.00   3500.00 1300.00      1
 1.09154411e+01 2.11069264e-02-1.04347901e-05 2.43633158e-09-2.20224945e-13    2
-1.35446352e+04-2.42468451e+01 1.81101363e+00 4.91205495e-02-4.27582013e-05    3
 1.90124399e-08-3.40793808e-12-1.11774841e+04 2.20654311e+01                   4
ZALD3OO                 C   3H   5O   5     G    300.00   3500.00 1800.00      1
 2.14549191e+01 1.08256409e-02-3.75393278e-06 5.88014012e-10-3.47282965e-14    2
-3.59900210e+04-7.93559882e+01 5.41191662e+00 4.64767576e-02-3.34631967e-05    3
 1.15914451e-08-1.56298261e-12-3.02145401e+04 7.47208817e+00                   4
ETC3H4O2                C   3H   4O   2     G    300.00   3500.00 1240.00      1
 1.02920429e+01 1.38871300e-02-6.12561993e-06 1.30548845e-09-1.09965765e-13    2
-3.57026988e+04-2.69350036e+01 1.17378044e-01 4.67086294e-02-4.58290467e-05    3
 2.26514168e-08-4.41358036e-12-3.31793820e+04 2.43405589e+01                   4
KEA3B3L                 C   3H   4O   4     G    300.00   3500.00 1500.00      1
 1.56495498e+01 1.47904716e-02-6.84032431e-06 1.49167146e-09-1.26830372e-13    2
-4.74213138e+04-4.92482738e+01 1.41905666e+00 5.27384532e-02-4.47883060e-05    3
 1.83574411e-08-2.93779198e-12-4.31521659e+04 2.51755980e+01                   4
RALD4OOX                C   4H   7O   3     G    300.00   3500.00 1060.00      1
 1.47280765e+01 1.68541717e-02-7.08657063e-07-1.32138238e-09 2.25378321e-13    2
-2.49490049e+04-4.17540781e+01-2.51677559e+00 8.19290853e-02-9.27957989e-05    3
 5.65950590e-08-1.34341597e-11-2.12930963e+04 4.24472035e+01                   4
QA4X                    C   4H   7O   3     G    300.00   3500.00 1020.00      1
 1.57879646e+01 1.38870673e-02 1.11593612e-06-1.77746725e-09 2.67503333e-13    2
-1.92489295e+04-4.33532546e+01-6.30635463e-01 7.82737344e-02-9.35703389e-05    3
 6.01089870e-08-1.49007453e-11-1.58995350e+04 3.61821314e+01                   4
ZA4X                    C   4H   7O   5     G    300.00   3500.00 1030.00      1
 2.21686912e+01 9.17757313e-03 7.13282539e-06-4.12053825e-09 5.56292343e-13    2
-3.97162883e+04-7.35383816e+01-2.33834122e+00 1.04350515e-01-1.31468546e-04    3
 8.55890871e-08-2.12178886e-11-3.46678396e+04 4.54182820e+01                   4
KEA4X                   C   4H   6O   4     G    300.00   3500.00  980.00      1
 1.51486382e+01 1.43075627e-02 4.47525531e-07-1.46947397e-09 2.26509070e-13    2
-1.74087245e+04-3.88103573e+01 7.77078059e-01 7.29669918e-02-8.93373148e-05    3
 5.96086487e-08-1.53546447e-11-1.45918987e+04 3.02337683e+01                   4
ETALD4X                 C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104167e+00 1.56985814e-02-7.47624893e-06 1.72107281e-09-1.55288692e-13    2
-3.54471815e+04-2.25395261e+01 7.88830836e-02 4.70057767e-02-4.66102431e-05    3
 2.34621807e-08-4.68468616e-12-3.31930634e+04 2.44846029e+01                   4
CH3COCHO                C   3H   4O   2     G    300.00   3500.00 1370.00      1
 1.06304440e+01 1.18394227e-02-4.21486308e-06 6.67473434e-10-3.88516159e-14    2
-4.37970340e+04-2.83088260e+01-8.46550190e-01 4.53488948e-02-4.09040660e-05    3
 1.85211002e-08-3.29681270e-12-4.06523375e+04 3.06741176e+01                   4
RALD5XOO                C   5H   9O   3     G    300.00   3500.00 1240.00      1
 5.00092606e+01-5.34134337e-02 6.46290203e-05-2.28767022e-08 2.64030383e-12    2
-4.06673538e+04-2.20829583e+02-1.12640294e+01 1.44242340e-01-1.74470706e-04    3
 1.05671538e-07-2.32766801e-11-2.54715779e+04 8.79592039e+01                   4
QA5X                    C   5H   9O   3     G    300.00   3500.00 1020.00      1
 3.16179276e+01-1.36493914e-02 3.39152688e-05-1.31900642e-08 1.56959131e-12    2
-3.26152700e+04-1.14322464e+02-3.56697746e+00 1.24330628e-01-1.68996525e-04    3
 1.19432023e-07-3.09358223e-11-2.54375494e+04 5.61211171e+01                   4
ZA5X                    C   5H   9O   5     G    300.00   3500.00 1030.00      1
 4.82844918e+01-4.15707481e-02 6.14657182e-05-2.30375148e-08 2.73823910e-12    2
-5.69207575e+04-1.98450742e+02-1.56034005e+01 2.06537571e-01-2.99857077e-04    3
 2.10828372e-07-5.40253257e-11-4.37598517e+04 1.11659857e+02                   4
KEA5X                   C   5H   8O   4     G    300.00   3500.00  890.00      1
 2.81159854e+01-1.51101029e-02 3.53666256e-05-1.35086149e-08 1.59169633e-12    2
 3.74972700e+04-9.42664385e+01 2.11579327e-01 1.10302958e-01-1.76003702e-04    3
 1.44821219e-07-4.28829760e-11 4.24642543e+04 3.71043837e+01                   4
RALD6XOO                C   6H  11O   3     G    300.00   3500.00 1240.00      1
 5.00092606e+01-5.34134337e-02 6.46290203e-05-2.28767022e-08 2.64030383e-12    2
-4.06673538e+04-2.20829583e+02-1.12640294e+01 1.44242340e-01-1.74470706e-04    3
 1.05671538e-07-2.32766801e-11-2.54715779e+04 8.79592039e+01                   4
QA6X                    C   6H  11O   3     G    300.00   3500.00 1020.00      1
 3.16179276e+01-1.36493914e-02 3.39152688e-05-1.31900642e-08 1.56959131e-12    2
-3.26152700e+04-1.14322464e+02-3.56697746e+00 1.24330628e-01-1.68996525e-04    3
 1.19432023e-07-3.09358223e-11-2.54375494e+04 5.61211171e+01                   4
ZA6X                    C   6H  11O   5     G    300.00   3500.00 1030.00      1
 4.82844918e+01-4.15707481e-02 6.14657182e-05-2.30375148e-08 2.73823910e-12    2
-5.69207575e+04-1.98450742e+02-1.56034005e+01 2.06537571e-01-2.99857077e-04    3
 2.10828372e-07-5.40253257e-11-4.37598517e+04 1.11659857e+02                   4
KEA6X                   C   6H  10O   4     G    300.00   3500.00  890.00      1
 2.81159854e+01-1.51101029e-02 3.53666256e-05-1.35086149e-08 1.59169633e-12    2
 3.74972700e+04-9.42664385e+01 2.11579328e-01 1.10302958e-01-1.76003702e-04    3
 1.44821219e-07-4.28829760e-11 4.24642543e+04 3.71043837e+01                   4
ETALD6X                 C   6H  10O   2     G    300.00   3500.00 1200.00      1
 9.47104167e+00 1.56985814e-02-7.47624893e-06 1.72107281e-09-1.55288692e-13    2
-3.54471815e+04-2.25395261e+01 7.88830836e-02 4.70057767e-02-4.66102431e-05    3
 2.34621807e-08-4.68468616e-12-3.31930634e+04 2.44846029e+01                   4
RIBALDGOO               C   4H   7O   3     G    300.00   3500.00 1090.00      1
 1.33433414e+01 1.84987671e-02-1.85145304e-06-9.50437233e-10 1.82631153e-13    2
-2.33799980e+04-3.43356040e+01-3.50808855e+00 8.03388770e-02-8.69525216e-05    3
 5.10991460e-08-1.17553467e-11-1.97063863e+04 4.84150219e+01                   4
RIBALDBOO               C   4H   7O   3     G    300.00   3500.00 1060.00      1
 1.47280765e+01 1.68541717e-02-7.08657063e-07-1.32138238e-09 2.25378321e-13    2
-2.49490049e+04-4.17540781e+01-2.51677559e+00 8.19290853e-02-9.27957989e-05    3
 5.65950590e-08-1.34341597e-11-2.12930963e+04 4.24472035e+01                   4
QIBALDG2                C   4H   7O   3     G    300.00   3500.00  980.00      1
 1.67965085e+01 1.08043172e-02 4.76341977e-06-3.20053120e-09 4.44231065e-13    2
-2.25755348e+04-5.02646403e+01-3.01325724e-01 8.05913956e-02-1.02053537e-04    3
 6.94640652e-08-1.80926558e-11-1.92243593e+04 3.18771037e+01                   4
QIBALDG3                C   4H   7O   3     G    300.00   3500.00 1050.00      1
 1.47854637e+01 1.55385624e-02-2.73488731e-07-1.29944016e-09 2.11492594e-13    2
-1.68282754e+04-3.82904661e+01-2.35309180e+00 8.08282978e-02-9.35445393e-05    3
 5.79202745e-08-1.38884395e-11-1.32291787e+04 4.52293503e+01                   4
QIBALDB3                C   4H   7O   3     G    300.00   3500.00 1020.00      1
 1.57879646e+01 1.38870673e-02 1.11593612e-06-1.77746725e-09 2.67503333e-13    2
-1.92489295e+04-4.33532546e+01-6.30635463e-01 7.82737344e-02-9.35703389e-05    3
 6.01089870e-08-1.49007453e-11-1.58995350e+04 3.61821314e+01                   4
ETIBALDGB               C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104167e+00 1.56985814e-02-7.47624893e-06 1.72107281e-09-1.55288692e-13    2
-3.54471815e+04-2.25395261e+01 7.88830836e-02 4.70057767e-02-4.66102431e-05    3
 2.34621807e-08-4.68468616e-12-3.31930634e+04 2.44846029e+01                   4
ETIBALDGG               C   4H   6O   2     G    300.00   3500.00 1200.00      1
 9.47104167e+00 1.56985814e-02-7.47624893e-06 1.72107281e-09-1.55288692e-13    2
-3.54471815e+04-2.25395261e+01 7.88830836e-02 4.70057767e-02-4.66102431e-05    3
 2.34621807e-08-4.68468616e-12-3.31930634e+04 2.44846029e+01                   4
ZIBALDG2                C   4H   7O   5     G    300.00   3500.00 1030.00      1
 2.21686912e+01 9.17757313e-03 7.13282539e-06-4.12053825e-09 5.56292343e-13    2
-3.97162883e+04-7.35383816e+01-2.33834122e+00 1.04350515e-01-1.31468546e-04    3
 8.55890871e-08-2.12178886e-11-3.46678396e+04 4.54182820e+01                   4
ZIBALDG3                C   4H   7O   5     G    300.00   3500.00 1080.00      1
 1.90668858e+01 1.53920232e-02 1.15889664e-06-1.93815091e-09 2.92451852e-13    2
-3.52242064e+04-5.68408680e+01-2.45362850e+00 9.50976318e-02-1.09543338e-04    3
 6.63965616e-08-1.55257686e-11-3.05757753e+04 4.86394149e+01                   4
ZIBALDB3                C   4H   7O   5     G    300.00   3500.00 1080.00      1
 1.90668858e+01 1.53920232e-02 1.15889664e-06-1.93815091e-09 2.92451852e-13    2
-3.52242064e+04-5.68408680e+01-2.45362850e+00 9.50976318e-02-1.09543338e-04    3
 6.63965616e-08-1.55257686e-11-3.05757753e+04 4.86394149e+01                   4
KIA4G2                  C   4H   6O   4     G    300.00   3500.00 1800.00      1
 2.35089845e+01 2.55786721e-03-1.96914845e-06 1.09436465e-09-1.65129977e-13    2
-5.44782542e+04-9.88855068e+01-1.84484588e+00 5.88997125e-02-4.89206862e-05    3
 1.84838231e-08-2.58033254e-12-4.53508752e+04 3.83347123e+01                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   3500.00 1470.00      1
 1.29296103e+01 3.16150611e-02-1.35584975e-05 2.81753187e-09-2.32686284e-13    2
-2.37933924e+04-4.88968549e+01-6.91462638e+00 8.56129840e-02-6.86584188e-05    3
 2.78061583e-08-4.48245269e-12-1.79591868e+04 5.44853543e+01                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   3500.00 1690.00      1
 2.24459936e+01 2.37621277e-02-8.83881474e-06 1.53830075e-09-1.04514815e-13    2
-5.03880249e+04-8.77405631e+01 1.27283562e+00 7.38761111e-02-5.33186817e-05    3
 1.90845993e-08-2.70012112e-12-4.32314975e+04 2.55178450e+01                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   3500.00 1660.00      1
 1.69989732e+01 3.01601499e-02-1.19254896e-05 2.25822367e-09-1.69878947e-13    2
-2.10464569e+04-6.14617731e+01 1.07910948e+00 6.85212672e-02-4.65891499e-05    3
 1.61793724e-08-2.26643749e-12-1.57610621e+04 2.34108339e+01                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   3500.00 1630.00      1
 1.86197530e+01 2.85111424e-02-1.13969334e-05 2.18137254e-09-1.65768942e-13    2
-1.50391446e+04-6.74883738e+01 1.48070310e+00 7.05701605e-02-5.01015514e-05    3
 1.80114821e-08-2.59369986e-12-9.45181437e+03 2.35714319e+01                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   3500.00 1800.00      1
 2.53088279e+01 2.46008468e-02-8.38584870e-06 1.28446216e-09-7.25492021e-14    2
-3.52662111e+04-9.88693150e+01 2.93992987e+00 7.43095092e-02-4.98097340e-05    3
 1.66266419e-08-2.20340750e-12-2.72134078e+04 2.21958278e+01                   4
CYC6-OO                 C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.87814621e+01 3.54361927e-02-1.49718784e-05 3.04328286e-09-2.46478319e-13    2
-1.95252830e+04-7.87240876e+01-6.50623568e+00 9.16310766e-02-6.18009483e-05    3
 2.03873828e-08-2.65538109e-12-1.04217118e+04 5.81382079e+01                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 1.91384147e+01 3.64873063e-02-1.63612962e-05 3.53264562e-09-3.02111689e-13    2
-1.43294351e+04-7.86383640e+01-4.87015408e+00 8.98396814e-02-6.08216088e-05    3
 1.99994281e-08-2.58916481e-12-5.68635037e+03 5.13010187e+01                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   3500.00 1800.00      1
 2.09300723e+01 3.28719793e-02-1.40160778e-05 2.89193638e-09-2.38539838e-13    2
-1.52994543e+04-8.89349636e+01-7.04914219e+00 9.50480115e-02-6.58294380e-05    3
 2.20820698e-08-2.90383614e-12-5.22693704e+03 6.24943819e+01                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.29323176e+01 2.20056554e-02-7.35242350e-06 1.07816406e-09-5.64635919e-14    2
-2.79806200e+04-1.10525203e+02-1.05629257e+01 9.64395294e-02-6.93806518e-05    3
 2.40515820e-08-3.24721608e-12-1.59223324e+04 7.07580407e+01                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.18028612e+01 2.41377428e-02-8.73118284e-06 1.46035609e-09-9.51866869e-14    2
-2.87387454e+04-1.06217525e+02-1.25990095e+01 1.00586344e-01-7.24383509e-05    3
 2.50556035e-08-3.37230438e-12-1.63540719e+04 7.99725758e+01                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   3500.00 1800.00      1
 2.14079592e+01 2.50825461e-02-9.38039634e-06 1.64525432e-09-1.14247640e-13    2
-3.89741817e+04-1.05728234e+02-1.45960517e+01 1.05091459e-01-7.60544907e-05    3
 2.63393633e-08-3.54398501e-12-2.60127378e+04 8.91329846e+01                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   3500.00 1800.00      1
 1.15965428e+01 4.02887933e-02-1.86685839e-05 4.15568433e-09-3.64030709e-13    2
-3.62221493e+04-4.27468435e+01-6.46490380e+00 8.04253413e-02-5.21157073e-05    3
 1.65435078e-08-2.08456175e-12-2.97200285e+04 5.50054734e+01                   4
C5H9CHO                 C   6H  10O   1     G    300.00   3500.00 1100.00      1
 9.07727161e+00 2.66919102e-02-7.89644695e-06 7.31227306e-10 1.61730960e-14    2
-1.68606427e+04-1.54909489e+01-3.32869064e-01 6.09106035e-02-5.45583015e-05    3
 2.90111392e-08-6.41107960e-12-1.47904117e+04 3.08044225e+01                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283790e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283790e-14    2
-3.55499047e+04-1.29752781e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.56593329e+01                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   3500.00 1770.00      1
 2.93742215e+01 2.67858800e-02-9.56345992e-06 1.54085681e-09-9.31283790e-14    2
-3.55499047e+04-1.30447295e+02-4.99061953e+00 1.04446538e-01-7.53775765e-05    3
 2.63296013e-08-3.59436348e-12-2.33847510e+04 5.49648189e+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.17655243e+01 3.67451403e-02-1.42717448e-05 2.74140448e-09-2.13135508e-13    2
-3.59903393e+04-5.10812501e+01-1.06696444e+01 9.82113560e-02-7.74219664e-05    3
 3.15771221e-08-5.15075839e-12-2.94392700e+04 6.56457555e+01                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415882e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.91587814e+01-8.02402159e+00 8.95009509e-02-6.86853397e-05    3
 2.77298319e-08-4.50893790e-12-3.06512867e+04 5.29538877e+01                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415882e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853397e-05    3
 2.77298319e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
C7DIONE                 C   7H  12O   2     G    300.00   3500.00  700.00      1
-7.55853626e-01 8.24536117e-02-4.58824666e-05 1.18274999e-08-1.15807940e-12    2
-3.67546789e+04 2.64722479e+01 3.52180416e+00 5.80098529e-02 6.49701649e-06    3
-3.80577221e-08 1.66580713e-11-3.73535510e+04 7.36075518e+00                   4
NC7H14O                 C   7H  14O   1     G    300.00   3500.00 1490.00      1
 1.37609323e+01 4.99379374e-02-2.21152348e-05 4.72010363e-09-3.98160015e-13    2
-3.97917916e+04-4.67908592e+01-7.39181742e+00 1.06723843e-01-7.92822536e-05    3
 3.02981881e-08-4.68978493e-12-3.34882722e+04 6.36941424e+01                   4
NC7H15-OO               C   7H  15O   2     G    300.00   3500.00 1780.00      1
 2.68006146e+01 3.35780867e-02-1.17982179e-05 1.89992230e-09-1.16218735e-13    2
-2.33388920e+04-1.06550436e+02 1.92333992e+00 8.94820746e-02-5.89083201e-05    3
 1.95441553e-08-2.59434135e-12-1.44825822e+04 2.78126029e+01                   4
NC7-QOOH                C   7H  15O   2     G    300.00   3500.00 1800.00      1
 3.67777501e+01 2.43465391e-02-1.65378816e-05 5.22869887e-09-5.85107382e-13    2
-2.84549794e+04-1.65059640e+02-2.87358792e+00 1.12460624e-01-8.99662853e-05    3
 3.24244039e-08-4.36228864e-12-1.41804977e+04 4.95416731e+01                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   3500.00 1690.00      1
 2.24694069e+01 4.29307086e-02-1.68910162e-05 3.18431082e-09-2.38592446e-13    2
-4.58962940e+04-7.93472401e+01 2.87430503e+00 8.93096479e-02-5.80557552e-05    3
 1.94228666e-08-2.64074567e-12-3.92731495e+04 2.54699082e+01                   4
C7KETONE                C   7H  14O   1     G    300.00   3500.00 1800.00      1
 1.82994273e+01 4.14393597e-02-1.71834162e-05 3.42714287e-09-2.72037363e-13    2
-4.27848802e+04-6.59785823e+01-2.29236271e-01 8.26141675e-02-5.14957561e-05    3
 1.61354169e-08-2.03707542e-12-3.61145614e+04 3.43024100e+01                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   3500.00 1670.00      1
 2.27584121e+01 4.25741258e-02-1.77950010e-05 3.55398723e-09-2.80791799e-13    2
-5.95329656e+04-8.19251638e+01 2.24997334e+00 9.16961348e-02-6.19165659e-05    3
 2.11673864e-08-2.91752820e-12-5.26831470e+04 2.75334100e+01                   4
NC7H15OOH               C   7H  16O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089265e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
IC8H16O                 C   8H  16O   1     G    300.00   3500.00 1730.00      1
 2.92525449e+01 3.42835226e-02-1.16024061e-05 1.77291875e-09-1.00401812e-13    2
-4.92824114e+04-1.33818841e+02-8.05235857e+00 1.20537635e-01-8.63892084e-05    3
 3.05924957e-08-4.26508057e-12-3.63749148e+04 6.66033697e+01                   4
IC8H17-OO               C   8H  17O   2     G    300.00   3500.00 1600.00      1
 2.43863221e+01 4.79091863e-02-1.96116165e-05 3.85759153e-09-3.01446048e-13    2
-3.51809040e+04-9.31491997e+01-7.10506923e-01 1.10651259e-01-7.84323095e-05    3
 2.83662136e-08-4.13091825e-12-2.71499187e+04 3.97240936e+01                   4
IC8-QOOH                C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574276e-02-1.91478836e-05 3.78861311e-09-2.97862013e-13    2
-2.91331926e+04-1.00455337e+02-9.92411233e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   3500.00 1560.00      1
 2.59202581e+01 4.65574276e-02-1.91478836e-05 3.78861311e-09-2.97862013e-13    2
-2.91331926e+04-1.00455337e+02-9.92411233e-01 1.15564272e-01-8.55006187e-05    3
 3.21444828e-08-4.84207190e-12-2.07364398e+04 4.13504180e+01                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   3500.00 1710.00      1
 3.48314225e+01 3.98146097e-02-1.43978345e-05 2.42273588e-09-1.57988116e-13    2
-5.01227380e+04-1.45334518e+02 1.76391327e+00 1.17165508e-01-8.22495001e-05    3
 2.88756269e-08-4.02536985e-12-3.88136498e+04 3.19375985e+01                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   3500.00 1770.00      1
 3.33140926e+01 3.48304479e-02-1.19632189e-05 1.85711682e-09-1.07309433e-13    2
-6.88276671e+04-1.40834098e+02 5.55148980e-01 1.08861959e-01-7.47017874e-05    3
 2.54874628e-08-3.44492892e-12-5.72310011e+04 3.59135548e+01                   4
KHDECA                  C  10H  16O   3     G    300.00   3500.00 1460.00      1
 1.16022418e+01 3.57303662e-02-1.34415882e-05 2.50437459e-09-1.89510289e-13    2
-3.63821557e+04-4.98532958e+01-8.02402159e+00 8.95009509e-02-6.86853397e-05    3
 2.77298319e-08-4.50893790e-12-3.06512867e+04 5.22593733e+01                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   3500.00 1650.00      1
 2.99089271e+01 5.87016385e-02-2.37959516e-05 4.63914803e-09-3.59659106e-13    2
-7.07246459e+04-1.14602343e+02 2.87865509e+00 1.24229571e-01-8.33667990e-05    3
 2.87081773e-08-4.00648172e-12-6.18046561e+04 2.93391873e+01                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762540e+01 8.51935060e-02-4.32222040e-05 1.03184896e-08-9.52873635e-13    2
-7.66784457e+04-1.07151303e+02 4.95723377e+00 1.38569107e-01-8.77018710e-05    3
 2.67924404e-08-3.24092235e-12-6.80315984e+04 2.28446447e+01                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1690.00      1
 4.88441297e+01 8.47833150e-02-3.17577492e-05 5.56702741e-09-3.82331486e-13    2
-9.50808904e+04-2.07202631e+02 1.75040693e+00 1.96247748e-01-1.30690678e-04    3
 4.45938236e-08-6.15552619e-12-7.91632121e+04 4.47087787e+01                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   3500.00 1590.00      1
 5.03105902e+01 8.85535013e-02-3.63077668e-05 7.13747183e-09-5.56692148e-13    2
-1.01978074e+05-2.30341253e+02-5.93668664e+00 2.30056085e-01-1.69800770e-04    3
 6.31093809e-08-9.35730677e-12-8.40914402e+04 6.71031189e+01                   4
IC12-OQOOH              C  12H  24O   3     G    300.00   3500.00 1800.00      1
 2.89762540e+01 8.51935060e-02-4.32222040e-05 1.03184896e-08-9.52873635e-13    2
-7.66784457e+04-1.07151303e+02 4.95723377e+00 1.38569107e-01-8.77018710e-05    3
 2.67924404e-08-3.24092235e-12-6.80315984e+04 2.28446447e+01                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.27624311e+01 3.77290665e-02-1.50512076e-05 2.88934934e-09-2.22140395e-13    2
-2.53740824e+04-9.90983226e+01-6.71698823e+00 1.03238887e-01-6.96427248e-05    3
 2.31084298e-08-3.03034602e-12-1.47614915e+04 6.04504445e+01                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522000e-06 1.12153176e-09-5.23348935e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   3500.00 1800.00      1
 2.93659891e+01 2.65374271e-02-8.30522000e-06 1.12153176e-09-5.23348935e-14    2
-2.28599204e+04-1.33867706e+02-7.82169678e+00 1.09176729e-01-7.71713049e-05    3
 2.66274891e-08-3.59482897e-12-9.47235352e+03 6.73998075e+01                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317082e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   3500.00 1770.00      1
 3.14587613e+01 3.12961497e-02-1.06604211e-05 1.62769455e-09-9.15073605e-14    2
-4.08526671e+04-1.40718316e+02-4.29317082e+00 1.12091476e-01-7.91310369e-05    3
 2.74170037e-08-3.73406515e-12-2.81964832e+04 5.21777121e+01                   4
KMCYC6                  C   7H  12O   3     G    300.00   3500.00 1800.00      1
 2.89245833e+01 2.89702632e-02-1.00807411e-05 1.60861341e-09-9.81376973e-14    2
-5.92858085e+04-1.29605491e+02-5.14358533e+00 1.04677305e-01-7.31699422e-05    3
 2.49749842e-08-3.34346697e-12-4.70212678e+04 5.47785441e+01                   4
QDECOOH                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
RDECOO                  C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
ZDECA                   C  10H  17O   4     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
DECA_ET                 C  10H  16O   1     G    300.00   3500.00 1450.00      1
 2.11071748e+01 5.53253918e-02-2.30739106e-05 4.67748686e-09-3.78388292e-13    2
-3.67326434e+04-9.38585120e+01-2.77500527e+01 1.90103951e-01-1.62500006e-04    3
 6.87814387e-08-1.14307938e-11-2.25640474e+04 1.60002934e+02                   4
NC10H21-OO              C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.23779830e+01 5.24885367e-02-1.93370131e-05 3.35369674e-09-2.28448799e-13    2
-4.06447276e+04-1.32098961e+02 1.67478189e+00 1.20717872e-01-7.61947929e-05    3
 2.44121337e-08-3.15323171e-12-2.95915752e+04 3.40731686e+01                   4
NC10-QOOH               C  10H  21O   2     G    300.00   3500.00 1800.00      1
 3.67714538e+01 4.56787199e-02-1.56929249e-05 2.49979255e-09-1.53467299e-13    2
-3.72897414e+04-1.54708984e+02 8.46533635e-01 1.25511876e-01-8.22205548e-05    3
 2.71396555e-08-3.57567048e-12-2.43567701e+04 3.97241784e+01                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   3500.00 1800.00      1
 4.08087722e+01 4.96339543e-02-1.81420129e-05 3.12006732e-09-2.11175643e-13    2
-5.65432959e+04-1.73811020e+02 2.62701325e+00 1.34482308e-01-8.88489740e-05    3
 2.93078307e-08-3.84836500e-12-4.27978627e+04 3.28366249e+01                   4
RODECOO                 C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
NC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763735e+01 5.51011625e-02-1.90602563e-05 3.05791504e-09-1.89217484e-13    2
-4.53973988e+04-1.84606456e+02 5.27389361e-01 1.49210016e-01-9.74843011e-05    3
 3.21038575e-08-4.22337617e-12-3.01517645e+04 4.45950809e+01                   4
NC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754174e+01 6.23046009e-02-2.29785783e-05 3.99220438e-09-2.72630412e-13    2
-4.86703034e+04-1.60846136e+02 1.39669302e+00 1.44257322e-01-9.12725124e-05    3
 2.92862540e-08-3.78569287e-12-3.53939626e+04 3.87492139e+01                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889668e+01 5.84439691e-02-2.09491581e-05 3.49897610e-09-2.27324947e-13    2
-6.45487872e+04-2.03262107e+02 2.75932352e+00 1.56509843e-01-1.02670720e-04    3
 3.37662211e-08-4.43110898e-12-4.86621157e+04 3.55767286e+01                   4
QODECOOH                C  10H  17O   2     G    300.00   3500.00 1800.00      1
 1.72379174e+01 3.76978745e-02-1.66331315e-05 3.54555182e-09-3.00284988e-13    2
-1.92027471e+04-7.01676462e+01-6.00367537e+00 8.93458584e-02-5.96731181e-05    3
 1.94862876e-08-2.51427606e-12-1.08357738e+04 5.56207021e+01                   4
IC12-QOOH               C  12H  25O   2     G    300.00   3500.00 1800.00      1
 4.28763735e+01 5.51011625e-02-1.90602563e-05 3.05791504e-09-1.89217484e-13    2
-4.53973988e+04-1.84606456e+02 5.27389361e-01 1.49210016e-01-9.74843011e-05    3
 3.21038575e-08-4.22337617e-12-3.01517645e+04 4.45950809e+01                   4
IC12H25-OO              C  12H  25O   2     G    300.00   3500.00 1800.00      1
 3.82754174e+01 6.23046009e-02-2.29785783e-05 3.99220438e-09-2.72630412e-13    2
-4.86703034e+04-1.60846136e+02 1.39669302e+00 1.44257322e-01-9.12725124e-05    3
 2.92862540e-08-3.78569287e-12-3.53939626e+04 3.87492139e+01                   4
IC12-OOQOOH             C  12H  25O   4     G    300.00   3500.00 1800.00      1
 4.68889668e+01 5.84439691e-02-2.09491581e-05 3.49897610e-09-2.27324947e-13    2
-6.45487872e+04-2.03262107e+02 2.75932352e+00 1.56509843e-01-1.02670720e-04    3
 3.37662211e-08-4.43110898e-12-4.86621157e+04 3.55767286e+01                   4
NC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.00344484e+01 8.20070153e-02-3.03042993e-05 5.28016700e-09-3.62022840e-13    2
-6.47045872e+04-2.18137205e+02 8.65096715e-01 1.91272241e-01-1.21358654e-04    3
 3.90040022e-08-5.04588884e-12-4.70036206e+04 4.79775838e+01                   4
IC16H33-OO              C  16H  33O   2     G    300.00   3500.00 1460.00      1
 3.94749769e+01 1.06211481e-01-4.74108472e-05 1.02029370e-08-8.67107397e-13    2
-6.81954459e+04-1.73182708e+02-7.55515778e+00 2.35061165e-01-1.79790660e-04    3
 7.06503399e-08-1.12176901e-11-5.44626465e+04 7.15084221e+01                   4
IC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1460.00      1
 4.22439745e+01 1.02589738e-01-4.54459634e-05 9.70909448e-09-8.19911244e-13    2
-6.26654622e+04-1.86283114e+02-7.79323360e+00 2.39677979e-01-1.86290047e-04    3
 7.40214614e-08-1.18323028e-11-4.80545975e+04 7.40533932e+01                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   3500.00 1560.00      1
 5.03537527e+01 8.72534729e-02-3.55849544e-05 6.99643634e-09-5.47405935e-13    2
-6.86134004e+04-2.32227161e+02-7.33743336e+00 2.35179591e-01-1.77821606e-04    3
 6.77813303e-08-1.02885748e-11-5.06137504e+04 7.17539151e+01                   4
NC16-QOOH               C  16H  33O   2     G    300.00   3500.00 1800.00      1
 5.49634696e+01 7.74662171e-02-2.71265902e-05 4.36953904e-09-2.68719606e-13    2
-8.49949222e+04-2.46825964e+02 8.02842617e-02 1.99428851e-01-1.28762119e-04    3
 4.20123273e-08-5.49688464e-12-6.52369755e+04 5.02132837e+01                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1800.00      1
 5.83925916e+01 7.87490302e-02-2.86987241e-05 4.90944001e-09-3.29403316e-13    2
-8.05061539e+04-2.59209019e+02 2.14519035e+00 2.03743255e-01-1.32860578e-04    3
 4.34879045e-08-5.68752339e-12-6.02570894e+04 4.52136503e+01                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   3500.00 1420.00      1
 4.21122112e+01 1.11834123e-01-5.11978482e-05 1.12541459e-08-9.72533984e-13    2
-7.89343498e+04-1.80495570e+02-6.54289827e+00 2.48890769e-01-1.95975996e-04    3
 7.92251073e-08-1.29392525e-11-6.51162987e+04 7.12984570e+01                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   3500.00 1370.00      1
 4.07769110e+01 1.15135971e-01-5.36319133e-05 1.19826916e-08-1.04989886e-12    2
-8.16821240e+04-1.74509322e+02-7.08781179e+00 2.54886986e-01-2.06643974e-04    3
 8.64411154e-08-1.46372025e-11-6.85671899e+04 7.14786263e+01                   4
RC6H5C4H8OO             C  10H  13O   2     G    300.00   3500.00 1800.00      1
 2.95255442e+01 3.88781010e-02-1.67600039e-05 3.28863590e-09-2.50060545e-13    2
-1.12745968e+04-1.27907262e+02-2.97080554e+00 1.11092212e-01-7.69384294e-05    3
 2.55769416e-08-3.34565856e-12 4.24089133e+02 4.79697618e+01                   4
QC6H5C4H8               C  10H  13O   2     G    300.00   3500.00 1600.00      1
 2.58642262e+01 4.31466453e-02-1.79342226e-05 3.56441659e-09-2.80425673e-13    2
-2.83088037e+03-1.02550382e+02-4.02896150e+00 1.17879615e-01-8.79963813e-05    3
 3.27569827e-08-4.84176413e-12 6.73493970e+03 5.57168755e+01                   4
QC6H5C4H8OO             C  10H  13O   4     G    300.00   3500.00 1340.00      1
 2.21297416e+01 5.89831670e-02-2.79882043e-05 6.34013620e-09-5.60973948e-13    2
-1.94753092e+04-7.75039096e+01-3.35040472e+00 1.35043305e-01-1.13130150e-04    3
 4.86993132e-08-8.46380548e-12-1.26466300e+04 5.28803321e+01                   4
KETBBZ                  C  10H  12O   3     G    300.00   3500.00 1370.00      1
 2.04509740e+01 5.51768971e-02-2.63137048e-05 5.98071386e-09-5.30329454e-13    2
-7.66936808e+03-7.18792904e+01-2.50633123e+00 1.22205525e-01-9.97027139e-05    3
 4.16931270e-08-7.04719318e-12-1.37906646e+03 4.61036429e+01                   4
NC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1800.00      1
 1.10496319e+01 1.81260731e-02-6.48607610e-06 1.10352513e-09-7.45033698e-14    2
-3.64580965e+04-3.27312856e+01-2.51644448e-01 4.32400205e-02-2.74143656e-05    3
 8.85474347e-09-1.15106147e-12-3.23896370e+04 2.84335795e+01                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 7.63374756e+00 2.08880310e-02-8.76974163e-06 1.80199756e-09-1.48384024e-13    2
-1.08851839e+04-1.05293244e+01 2.18301336e+00 3.30007737e-02-1.88636939e-05    3
 5.54049839e-09-6.67620249e-13-8.92291955e+03 1.89711862e+01                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.06992300e+01 1.62004106e-02-6.03307514e-06 1.08996004e-09-7.93898637e-14    2
-1.44167384e+04-2.94436050e+01 9.48802516e-01 3.78680272e-02-2.40894223e-05    3
 7.77749601e-09-1.00821430e-12-1.09065845e+04 2.33277424e+01                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   3500.00 1800.00      1
 1.10024651e+01 1.50905454e-02-5.07771786e-06 7.82747262e-10-4.56159151e-14    2
-1.15495011e+04-2.90815232e+01 2.77594410e-01 3.89235914e-02-2.49385895e-05    3
 8.13862564e-09-1.06726569e-12-7.68854770e+03 2.89637142e+01                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   3500.00 1800.00      1
 6.66433268e+00 2.45624525e-02-1.14187516e-05 2.58003280e-09-2.29895788e-13    2
-7.91390086e+03-8.44862881e+00 1.62185706e+00 3.57679539e-02-2.07566695e-05    3
 6.03852088e-09-7.10241355e-13-6.09860964e+03 1.88423012e+01                   4
IC3H7OH                 C   3H   8O   1     G    300.00   3500.00 1490.00      1
 1.02736687e+01 1.89903342e-02-6.50928762e-06 9.85863990e-10-5.35101895e-14    2
-3.77812744e+04-2.92304676e+01-1.25951086e+00 4.99518902e-02-3.76786393e-05    3
 1.49318826e-08-2.39344620e-12-3.43443869e+04 3.10096138e+01                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   3500.00 1380.00      1
 6.32694430e+00 2.38762490e-02-1.07376178e-05 2.33737032e-09-2.01069469e-13    2
-1.14217376e+04-3.95690498e+00 6.40756936e-01 4.03579515e-02-2.86525118e-05    3
 1.09919085e-08-1.76892059e-12-9.85234986e+03 2.53070892e+01                   4
CH3COHCH3               C   3H   7O   1     G    300.00   3500.00 1270.00      1
 6.71652579e+00 2.35306498e-02-1.06144747e-05 2.31761627e-09-1.99886320e-13    2
-1.44175086e+04-7.90476331e+00 1.21649821e+00 4.08535713e-02-3.10746182e-05    3
 1.30578491e-08-2.31410538e-12-1.30205016e+04 1.99442900e+01                   4
C3H7CHO                 C   4H   8O   1     G    300.00   3500.00  700.00      1
-9.77279407e-01 5.24983746e-02-3.09762337e-05 8.32680249e-09-8.38156518e-13    2
-2.70767712e+04 3.27194911e+01 3.71554479e+00 2.56822364e-02 2.64869197e-05    3
-4.64000103e-08 1.87071338e-11-2.77337665e+04 1.17531399e+01                   4
RALD4X                  C   4H   7O   1     G    300.00   3500.00 1140.00      1
-3.84911251e+00 5.11968669e-02-2.73583537e-05 6.64027831e-09-6.13455715e-13    2
-5.69209146e+03 4.92440537e+01 6.06312506e+00 1.64170860e-02 1.84045160e-05    3
-2.01216338e-08 5.25538465e-12-7.95208163e+03 1.24454033e-01                   4
C3H5CHO                 C   4H   6O   1     G    300.00   3500.00 1610.00      1
 9.36564259e+00 1.99394689e-02-8.24714277e-06 1.63840913e-09-1.29181894e-13    2
-1.44293663e+04-2.07054000e+01 2.40474771e-01 4.26106933e-02-2.93694015e-05    3
 1.03846860e-08-1.48729943e-12-1.14910622e+04 2.76639767e+01                   4
IC3H5CHO                C   4H   6O   1     G    300.00   3500.00 1370.00      1
 8.96605760e+00 2.20962385e-02-1.00901145e-05 2.22139279e-09-1.91792264e-13    2
-1.79920102e+04-2.11939239e+01 6.92941976e-01 4.62513206e-02-3.65372847e-05    3
 1.50910620e-08-2.54027204e-12-1.57251765e+04 2.13235423e+01                   4
NC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1260.00      1
 9.47752943e+00 2.59932961e-02-1.14395843e-05 2.45196196e-09-2.08596763e-13    2
-2.58308658e+04-2.26233180e+01-1.20059161e+00 5.98920930e-02-5.17952949e-05    3
 2.38041898e-08-4.44514991e-12-2.31399793e+04 3.13602824e+01                   4
IC4H7OH                 C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.15391986e+01 2.16392182e-02-8.55965721e-06 1.65851647e-09-1.29717162e-13    2
-2.50645509e+04-3.36074037e+01 1.41746535e+00 4.41319587e-02-2.73036076e-05    3
 8.60072033e-09-1.09391214e-12-2.14207270e+04 2.11735281e+01                   4
IC3H7CHO                C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.25375038e+01 2.06759832e-02-7.90606663e-06 1.44761601e-09-1.05776578e-13    2
-3.22363635e+04-4.10505202e+01-3.44732114e-01 4.93031741e-02-3.17620591e-05    3
 1.02831688e-08-1.33293668e-12-2.75987585e+04 2.86708279e+01                   4
RIBALDB                 C   4H   7O   1     G    300.00   3500.00 1090.00      1
 7.80130143e+00 2.08311674e-02-4.31906593e-06-1.13870083e-10 8.81387266e-14    2
-1.58031223e+03-1.28298252e+01-1.99174484e+00 5.67689519e-02-5.37747327e-05    3
 3.01342441e-08-6.84950215e-12 5.54571859e+02 3.52599043e+01                   4
RIBALDG                 C   4H   7O   1     G    300.00   3500.00 1050.00      1
 9.00440173e+00 1.88029635e-02-3.43463806e-06-2.58096325e-10 9.53220855e-14    2
-4.96767967e+03-1.61872934e+01-3.42297331e+00 6.61453446e-02-7.10666111e-05    3
 4.26828389e-08-1.01287101e-11-2.35793091e+03 4.43739411e+01                   4
N1C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.48230798e+01 2.16832754e-02-7.46704085e-06 1.19388940e-09-7.36745676e-14    2
-4.08306213e+04-5.15940698e+01-4.78997489e-01 5.56878916e-02-3.58042210e-05    3
 1.16891413e-08-1.53134844e-12-3.53218735e+04 3.12239645e+01                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.13530982e+01 2.45578872e-02-9.82948618e-06 1.91527532e-09-1.49940483e-13    2
-1.52382167e+04-2.90980437e+01 1.95582522e+00 4.54407161e-02-2.72318436e-05    3
 8.36059288e-09-1.04512348e-12-1.18551985e+04 2.17619582e+01                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   3500.00 1790.00      1
 1.44669850e+01 1.91857603e-02-6.39892959e-06 9.65852776e-10-5.40086293e-14    2
-1.57844512e+04-4.62017057e+01 4.01250150e-02 5.14245536e-02-3.34146782e-05    3
 1.10275841e-08-1.45927837e-12-1.06196353e+04 3.17990977e+01                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 9.76394270e+00 2.97115921e-02-1.36105451e-05 3.01462692e-09-2.63554924e-13    2
-1.20864790e+04-2.37714276e+01 1.13482603e+00 4.88874069e-02-2.95903908e-05    3
 8.93308828e-09-1.08556345e-12-8.97999699e+03 2.29311520e+01                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.45806677e+01 1.95400847e-02-6.85981976e-06 1.13500508e-09-7.38190524e-14    2
-1.88304378e+04-4.88995705e+01 7.07705507e-01 5.03688897e-02-3.25504906e-05    3
 1.06500683e-08-1.39535562e-12-1.38361714e+04 2.61837951e+01                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.10474004e+01 2.49495870e-02-1.02454957e-05 2.07975625e-09-1.70767943e-13    2
-1.60937900e+04-2.75546799e+01-8.85955889e-02 4.96962447e-02-3.08677104e-05    3
 9.71761356e-09-1.23158146e-12-1.20848314e+04 3.27156533e+01                   4
N2C4H9OH                C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.39850075e+01 2.35768220e-02-8.73106105e-06 1.51546162e-09-1.02847459e-13    2
-4.24053999e+04-4.83702850e+01 1.11912947e-01 5.44059211e-02-3.44219770e-05    3
 1.10306157e-08-1.42439663e-12-3.74110858e+04 2.67137971e+01                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097164e-06 1.27900113e-09-8.37238499e-14    2
-1.74897435e+04-4.46134901e+01 9.11733055e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.39333095e+01 2.07599768e-02-7.56097164e-06 1.27900113e-09-8.37238499e-14    2
-1.74897435e+04-4.46134901e+01 9.11733055e-01 4.96968134e-02-3.16750021e-05    3
 1.02101235e-08-1.32415752e-12-1.28019760e+04 2.58619981e+01                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   3500.00 1800.00      1
 1.11524016e+01 2.52912378e-02-1.05179486e-05 2.12392651e-09-1.71553011e-13    2
-1.78095410e+04-2.94209720e+01 6.76902372e-01 4.85701251e-02-2.99170213e-05    3
 9.30876824e-09-1.16944770e-12-1.40383613e+04 2.72746153e+01                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   3500.00 1430.00      1
 8.72382272e+00 3.04342830e-02-1.39185549e-05 3.06043861e-09-2.64689230e-13    2
-1.80661273e+04-1.71435098e+01 1.27395834e+00 5.12730645e-02-3.57774166e-05    3
 1.32510501e-08-2.04626467e-12-1.59354661e+04 2.14624055e+01                   4
TC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1440.00      1
 9.08150387e+00 3.22201837e-02-1.41979352e-05 3.03249263e-09-2.56658356e-13    2
-4.23917231e+04-2.36263218e+01-6.99999563e-01 5.93910266e-02-4.25008966e-05    3
 1.61357155e-08-2.53152343e-12-3.95746501e+04 2.71305359e+01                   4
RTC4H8OH                C   4H   9O   1     G    300.00   3500.00 1380.00      1
 8.66823484e+00 3.01271731e-02-1.35256253e-05 2.94117291e-09-2.52822189e-13    2
-1.73478965e+04-1.68023720e+01 1.39901310e-03 5.52484364e-02-4.08313463e-05    3
 1.61323424e-08-2.64252681e-12-1.49558499e+04 2.78015457e+01                   4
IC4H9OH                 C   4H  10O   1     G    300.00   3500.00 1800.00      1
 1.44537517e+01 2.20810695e-02-7.57959310e-06 1.19533670e-09-7.16167606e-14    2
-4.15822810e+04-5.13315495e+01-5.45479447e-01 5.54126942e-02-3.53559470e-05    3
 1.14828752e-08-1.50044155e-12-3.61825578e+04 2.98474183e+01                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   3500.00 1450.00      1
 8.91411879e+00 2.94184843e-02-1.30488503e-05 2.81020956e-09-2.39749810e-13    2
-1.71145335e+04-1.85255698e+01 6.16106328e-01 5.23095531e-02-3.67292664e-05    3
 1.36977572e-08-2.11691319e-12-1.47081099e+04 2.45907827e+01                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   3500.00  700.00      1
 2.02076660e+00 4.09903684e-02-2.06486867e-05 5.00507650e-09-4.71523454e-13    2
-1.40718373e+04 2.15880988e+01 3.53447956e+00 3.23405800e-02-2.11342588e-06    3
-1.26475529e-08 5.83298703e-12-1.42837571e+04 1.48252122e+01                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   3500.00 1780.00      1
 1.38129919e+01 2.02819032e-02-7.03372780e-06 1.12439860e-09-6.86002895e-14    2
-1.64045579e+04-4.42517079e+01 2.32452600e-01 5.07999690e-02-3.27511989e-05    3
 1.07564103e-08-1.42141092e-12-1.15698860e+04 2.90972641e+01                   4
MEK                     C   4H   8O   1     G    300.00   3500.00 1800.00      1
 1.00996674e+01 2.22850926e-02-8.24112797e-06 1.42760366e-09-9.77654879e-14    2
-3.40270944e+04-2.55002808e+01 1.67138626e+00 4.10146063e-02-2.38490560e-05    3
 7.20831776e-09-9.00642447e-13-3.09929132e+04 2.01153350e+01                   4
C5H9OH                  C   5H  10O   1     G    300.00   3500.00 1210.00      1
 1.31847853e+01 3.05720306e-02-1.32292735e-05 2.77400243e-09-2.30719149e-13    2
-2.99739271e+04-4.19054228e+01-3.87325759e+00 8.69622549e-02-8.31345102e-05    3
 4.12892844e-08-8.18842203e-12-2.58458807e+04 4.36413837e+01                   4
C4H9CHO                 C   5H  10O   1     G    300.00   3500.00  760.00      1
-1.78433184e+00 6.31204388e-02-3.60836199e-05 9.48321924e-09-9.39522549e-13    2
-2.97113508e+04 3.92478714e+01 5.53299033e+00 2.46082168e-02 3.99273445e-05    3
-5.71930654e-08 2.09934658e-11-3.08235838e+04 5.95416457e+00                   4
IC5H9OH                 C   5H  10O   1     G    300.00   3500.00 1340.00      1
 1.04339676e+01 3.43709884e-02-1.53823526e-05 3.33540372e-09-2.86051918e-13    2
-3.01866098e+04-2.68956309e+01-1.89607142e+00 7.11770751e-02-5.65831958e-05    3
 2.38333357e-08-4.11029295e-12-2.68821593e+04 3.61983077e+01                   4
IC4H9CHO                C   5H  10O   1     G    300.00   3500.00 1800.00      1
 1.47934378e+01 2.65660103e-02-1.04284281e-05 1.98344196e-09-1.51387846e-13    2
-3.60342983e+04-5.12505581e+01 7.73443177e-01 5.77215539e-02-3.63913811e-05    3
 1.15993505e-08-1.48693069e-12-3.09871002e+04 2.46285774e+01                   4
RALD5X                  C   5H   9O   1     G    300.00   3500.00  750.00      1
-3.04813122e-01 5.67977503e-02-3.24057644e-05 8.50471990e-09-8.41763295e-13    2
-5.21420509e+03 3.41933262e+01 6.22525357e+00 2.19707280e-02 3.72482804e-05    3
-5.34099865e-08 1.97964722e-11-6.19371509e+03 4.56811230e+00                   4
ALDC6                   C   6H  12O   1     G    300.00   3500.00 1800.00      1
 1.43376050e+01 3.78182965e-02-1.64821906e-05 3.50929997e-09-2.98005833e-13    2
-3.75955824e+04-4.53859600e+01 1.31726275e+00 6.67523904e-02-4.05939354e-05    3
 1.24395759e-08-1.53832193e-12-3.29082592e+04 2.50828483e+01                   4
RALD6X                  C   6H  11O   1     G    300.00   3500.00 1160.00      1
 5.47459470e-01 6.16901246e-02-2.98352974e-05 6.64392083e-09-5.73135815e-13    2
-1.27523068e+04 2.98980226e+01 4.05975345e+00 4.95787661e-02-1.41740579e-05    3
-2.35679152e-09 1.36667288e-12-1.35671590e+04 1.24319397e+01                   4
C5H11OH                 C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.84921366e+01 2.54355952e-02-8.57802272e-06 1.32118635e-09-7.66433346e-14    2
-4.51605186e+04-6.98750288e+01-6.77485013e-01 6.80347542e-02-4.40773219e-05    3
 1.44690750e-08-1.90273897e-12-3.82594548e+04 3.38749622e+01                   4
RPENT1OHA               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.84065773e+01 2.29900185e-02-7.76357329e-06 1.20244128e-09-7.05741185e-14    2
-2.32226149e+04-6.80495353e+01 4.75636951e-01 6.28365526e-02-4.09690184e-05    3
 1.35007543e-08-1.77867315e-12-1.67674764e+04 2.89964546e+01                   4
RPENT1OHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.50707231e+01 2.82315427e-02-1.08918053e-05 2.02927093e-09-1.51568857e-13    2
-1.95906718e+04-4.76575366e+01 1.72826109e+00 5.78814583e-02-3.56000684e-05    3
 1.11804795e-08-1.42257004e-12-1.47873854e+04 2.45546514e+01                   4
IC5H11OH                C   5H  12O   1     G    300.00   3500.00 1800.00      1
 1.75261800e+01 2.67328515e-02-9.21962742e-06 1.46158882e-09-8.81568439e-14    2
-4.58408793e+04-6.62686894e+01-6.91392019e-01 6.72163448e-02-4.29558718e-05    3
 1.39564942e-08-1.82356036e-12-3.92825534e+04 3.23286106e+01                   4
RIPENTOHA               C   5H  11O   1     G    300.00   3500.00 1620.00      1
 1.36179105e+01 3.09491059e-02-1.25439310e-05 2.45214936e-09-1.90908871e-13    2
-2.20274849e+04-4.25086987e+01 6.58084780e-01 6.29486755e-02-4.21731621e-05    3
 1.46452486e-08-2.07255998e-12-1.78285014e+04 2.62671274e+01                   4
RIPENTOHB               C   5H  11O   1     G    300.00   3500.00 1800.00      1
 1.43827445e+01 2.99341363e-02-1.24371812e-05 2.55513031e-09-2.11814101e-13    2
-2.12442482e+04-4.60019499e+01-6.44588846e-01 6.33282104e-02-4.02655763e-05    3
 1.28619433e-08-1.64331591e-12-1.58344082e+04 3.53291130e+01                   4
C6H13OH                 C   6H  14O   1     G    300.00   3500.00 1800.00      1
 2.78613474e+01 1.77437818e-02-2.99502852e-06 1.18974668e-11 2.84572872e-14    2
-5.19282550e+04-1.19896980e+02-1.83303781e+00 8.37313045e-02-5.79846308e-05    3
 2.03784168e-08-2.80022596e-12-4.12382763e+04 4.08152273e+01                   4
RHEX1OHA                C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.84298178e+01 1.33218304e-02-9.68178066e-07-3.32583082e-10 4.90833295e-14    2
-3.02913834e+04-1.20327849e+02-1.87679570e-01 7.69162690e-02-5.39635435e-05    3
 1.92953301e-08-2.67701572e-12-1.99890844e+04 3.45560167e+01                   4
RHEX1OHB                C   6H  13O   1     G    300.00   3500.00 1800.00      1
 2.97416428e+01 1.08284395e-02 6.26458140e-07-7.76125692e-10 9.43842404e-14    2
-2.87904782e+04-1.27477419e+02-8.09485399e-02 7.71008646e-02-5.46005628e-05    3
 1.96783265e-08-2.74651190e-12-1.80543453e+04 3.39286664e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559082e+01 1.49866375e-02-1.56738310e-06-4.84518439e-10 9.00436513e-14    2
-2.80668702e+04-9.05497671e+01-1.97000865e+00 6.65997861e-02-4.45783403e-05    3
 1.54454657e-08-2.12245414e-12-1.97055401e+04 3.51537401e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93193785e+00 3.75440987e-02-1.65478566e-05 3.53633643e-09-2.99976701e-13    2
-1.73087074e+03-8.88710671e+00-3.57520449e+00 6.08933039e-02-3.60055276e-05    3
 1.07428812e-08-1.30088570e-12 2.05170050e+03 4.79797395e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220811e+01 2.73824077e-02-1.01392581e-05 1.77707009e-09-1.22756971e-13    2
-2.85197010e+04-6.62488521e+01-2.62463459e+00 7.07864445e-02-4.84369376e-05    3
 1.67957680e-08-2.33138901e-12-2.22478177e+04 3.25342362e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276289e+01 2.66845577e-02-1.02158264e-05 1.86929104e-09-1.35803312e-13    2
-2.94216421e+03-5.15145769e+01-1.29689709e+00 6.41085720e-02-4.38302105e-05    3
 1.52882069e-08-2.14462305e-12 2.27642747e+03 3.18773552e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929736e+01 2.82582223e-02-1.13863841e-05 2.22526491e-09-1.74280993e-13    2
-1.02483443e+04-3.39253533e+01-6.89551965e-01 5.46638348e-02-3.33910611e-05    3
 1.03751453e-08-1.30620882e-12-5.97063504e+03 3.03853541e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
B1M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.21299340e+01 2.65376145e-02-1.02995525e-05 1.93064538e-09-1.45051208e-13    2
-1.11266091e+04-3.96207198e+01-6.39002025e-01 5.49130280e-02-3.39457304e-05    3
 1.06884890e-08-1.36141838e-12-6.52979211e+03 2.94874259e+01                   4
B1M3                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.31681365e+01 2.49963287e-02-9.30063098e-06 1.64277853e-09-1.14892348e-13    2
-1.09953810e+04-4.60629131e+01-8.44094903e-01 5.61346208e-02-3.52492077e-05    3
 1.12533625e-08-1.44969568e-12-5.95097767e+03 2.97742066e+01                   4
B2M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 9.73411699e+00 3.08235227e-02-1.30972997e-05 2.71635425e-09-2.25270435e-13    2
-1.14704814e+04-2.74877025e+01 1.14407401e-01 5.22006552e-02-3.09115767e-05    3
 9.31423462e-09-1.14164271e-12-8.00738598e+03 2.45761726e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099916e+00 2.71082714e-02-1.07932861e-05 1.95387665e-09-1.31111174e-13    2
-1.09862538e+03-2.37608448e+01-6.56863981e+00 6.82031726e-02-5.30140751e-05    3
 2.12327757e-08-3.43229252e-12 3.28126920e+03 5.42801525e+01                   4
LC5H8                   C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829160e+00 2.51033002e-02-8.43679233e-06 8.19905618e-10 3.11426514e-14    2
 4.67953300e+03-2.40439629e+01 1.19183501e+00 4.68276543e-02-3.12245763e-05    3
 1.14435811e-08-1.82614328e-12 6.90073958e+03 1.62025638e+01                   4
CYC5H7                  C   5H   7          G    200.00   3500.00 1740.00      1
 1.46691728e+01 1.34698305e-02-2.95655819e-06 2.78903446e-11 3.93991651e-14    2
 1.32998383e+04-5.70832491e+01-3.51544371e+00 5.52735467e-02-3.89942446e-05    3
 1.38354330e-08-1.94444317e-12 1.96280848e+04 4.07192024e+01                   4
LC5H7                   C   5H   7          G    200.00   3500.00 1640.00      1
 1.25568519e+01 1.79546663e-02-5.75033141e-06 7.12773055e-10-2.19484675e-14    2
 1.85872287e+04-4.12604534e+01-8.15591381e-01 5.05703817e-02-3.55817784e-05    3
 1.28393775e-08-1.87051622e-12 2.29733901e+04 2.98691530e+01                   4
DIALLYL                 C   6H  10          G    300.00   3500.00 1670.00      1
 1.46885479e+01 2.58341295e-02-9.34005191e-06 1.60362032e-09-1.08722036e-13    2
 2.72208305e+03-5.11904321e+01-8.93391062e-01 6.31561390e-02-4.28628150e-05    3
 1.49859609e-08-2.11206643e-12 7.92645066e+03 3.19742028e+01                   4
RC6H9A                  C   6H   9          G    300.00   3500.00 1310.00      1
 1.02179198e+01 3.31131696e-02-1.50182300e-05 3.28859653e-09-2.83959224e-13    2
 2.30740211e+04-2.53806643e+01-2.61882183e+00 7.23093274e-02-5.98993266e-05    3
 2.61288493e-08-4.64278609e-12 2.64372474e+04 4.00154625e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772261e+00 3.45074855e-02-1.63846780e-05 3.69260974e-09-3.24421025e-13    2
 5.74022138e+03-2.73566208e+01-6.91358136e+00 7.63364895e-02-5.84944135e-05    3
 2.25336547e-08-3.48567018e-12 1.03834500e+04 5.40276160e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624858e+01 2.76360017e-02-1.05259858e-05 1.89586361e-09-1.35054774e-13    2
-9.29985244e+03-6.25064559e+01-6.01517655e+00 7.46974737e-02-4.97438791e-05    3
 1.64210093e-08-2.15243611e-12-1.67589399e+03 5.21114707e+01                   4
RCYC6H9                 C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670463e+01 2.75651338e-02-1.13337615e-05 2.23021652e-09-1.74683445e-13    2
 7.93866332e+03-5.85441979e+01-6.48639356e+00 7.34616669e-02-4.95808724e-05    3
 1.63958131e-08-2.14212742e-12 1.53739017e+04 5.32365273e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578097e+01 4.34354098e-02-2.02455774e-05 4.54245292e-09-4.01195170e-13    2
-2.30439963e+04-4.47863376e+01-9.43363126e+00 8.94163897e-02-5.85630607e-05    3
 1.87341134e-08-2.37225913e-12-1.55950776e+04 6.72000574e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879191e+01 3.94798364e-02-1.80474738e-05 3.97976998e-09-3.47933572e-13    2
 4.69934404e+02-4.15743644e+01-9.20200373e+00 8.50129981e-02-5.59917752e-05    3
 1.80332150e-08-2.29980093e-12 7.84630661e+03 6.93213721e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951655e+01 5.24635940e-03 6.43208140e-06-3.19131390e-09 4.01093698e-13    2
-1.79767847e+04-1.24497292e+02-1.85358315e+00 7.25469181e-02-5.02818725e-05    3
 1.80498674e-08-2.58221828e-12-7.31503024e+03 3.72569567e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696120e+01 1.73458864e-02-4.57663866e-07-1.06280964e-09 1.59098857e-13    2
-3.76541592e+04-1.40920498e+02-2.76912812e+00 9.25430866e-02-6.31219974e-05    3
 2.21462028e-08-3.06437509e-12-2.54722127e+04 4.22218230e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938298e+01 4.32851195e-02-1.83429598e-05 3.81524631e-09-3.18291961e-13    2
-8.33589206e+03-5.34387877e+01-1.03213606e+00 8.08983770e-02-4.96873411e-05    3
 1.54242764e-08-1.93065725e-12-2.24254435e+03 3.81680706e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668105e+01 3.59607889e-02-1.37346402e-05 2.52229049e-09-1.85248240e-13    2
-1.87497345e+04-6.92309266e+01-1.22797310e+00 7.92825302e-02-4.98360912e-05    3
 1.58931983e-08-2.04231877e-12-1.17316124e+04 3.62789089e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155885e+01 4.43694094e-02-1.35968858e-05 1.75327621e-09-6.83090867e-14    2
-3.76580614e+04-8.42148794e+01-5.96912082e+00 1.20872170e-01-9.61538218e-05    3
 4.13489290e-08-7.18982937e-12-3.02675122e+04 5.27954202e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104230e+01 3.01796816e-02-5.82184988e-06 1.42085775e-11 7.60110768e-14    2
-1.80373025e+04-1.14981197e+02-3.32961207e+00 1.08192845e-01-8.23053436e-05    3
 3.33403496e-08-5.36943681e-12-8.90625182e+03 4.16697270e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616063e+01 4.14292819e-02-1.28170543e-05 1.66806735e-09-6.58961701e-14    2
-2.24684067e+04-7.38514297e+01-5.35586582e+00 1.10622059e-01-8.69521730e-05    3
 3.69705048e-08-6.36990286e-12-1.56875145e+04 5.11323812e+01                   4
DIMEPTD                 C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755546e+01 3.27318282e-02-1.05955708e-05 1.52102629e-09-7.69415904e-14    2
-6.19682930e+03-5.37226047e+01-1.29247814e+00 8.36265847e-02-6.88720095e-05    3
 3.11782470e-08-5.73671653e-12-1.82980473e+03 3.11918394e+01                   4
C7H8                    C   7H   8          G    200.00   3500.00 1740.00      1
 1.92535108e+01 1.64137602e-02-3.61135948e-06 2.27424890e-11 5.04456794e-14    2
-3.67626229e+03-8.27561068e+01-4.42382865e+00 7.08444256e-02-5.05343469e-05    3
 1.80008986e-08-2.53262272e-12 4.56345183e+03 4.45878951e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867713e+01 2.02277643e-02-7.36599497e-06 1.21196287e-09-7.46105009e-14    2
-1.80542263e+04-5.08485812e+01-5.47325436e+00 7.87541571e-02-7.33732049e-05    3
 3.42982837e-08-6.29384373e-12-1.28778595e+04 4.85843830e+01                   4
C6H5CHO                 C   7H   6O   1     G    200.00   3500.00 1630.00      1
 2.06104936e+01 1.34209230e-02-2.83635978e-06-5.48103780e-11 5.23167108e-14    2
-1.43315560e+04-8.70895599e+01-3.50845143e+00 7.26085180e-02-5.73034718e-05    3
 2.22221271e-08-3.36439149e-12-6.46877992e+03 4.10544422e+01                   4
C6H5CO                  C   7H   5O   1     G    300.00   3500.00 1470.00      1
 1.31799087e+01 2.42895707e-02-1.09067387e-05 2.35371847e-09-2.00195165e-13    2
 5.86598787e+03-4.37756649e+01-1.56203256e+00 6.44036967e-02-5.18395203e-05    3
 2.09173383e-08-3.35727336e-12 1.02001186e+04 3.30251959e+01                   4
C7H7                    C   7H   7          G    200.00   3500.00 1600.00      1
 1.77148781e+01 1.72901839e-02-4.74309316e-06 3.88421745e-10 1.27959347e-14    2
 1.68881058e+04-7.24712964e+01-3.23806381e+00 6.96725387e-02-5.38515508e-05    3
 2.08502791e-08-3.18436927e-12 2.35930472e+04 3.84624951e+01                   4
CH3C6H4                 C   7H   7          G    200.00   3500.00 1730.00      1
 1.83842182e+01 1.52647348e-02-3.43004339e-06 5.73661650e-11 4.21798063e-14    2
 2.84624024e+04-7.44700925e+01-2.82564598e+00 6.43048832e-02-4.59504033e-05    3
 1.64428613e-08-2.32566631e-12 3.58010154e+04 3.94808224e+01                   4
C6H5O                   H   5C   6O   1     G    100.00   3500.00 1800.00      1
 1.20320192e+01 2.29423311e-02-1.10171059e-05 2.53057377e-09-2.25735901e-13    2
 2.17286268e+02-4.10084349e+01 4.06305309e-01 4.87772509e-02-3.25462057e-05    3
 1.05043144e-08-1.33319988e-12 4.40254327e+03 2.19123540e+01                   4
CYC6H4                  C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465819e+01 1.50373245e-02-5.27844957e-06 8.14607575e-10-4.49073360e-14    2
 5.03301418e+04-3.53782935e+01-3.73796174e+00 5.69931634e-02-5.02311341e-05    3
 2.22206478e-08-3.86741452e-12 5.44418140e+04 4.04070822e+01                   4
OC6H4OH                 H   5C   6O   2     G    200.00   3500.00 1330.00      1
 9.78515606e+00 3.14205686e-02-1.61320626e-05 4.01581601e-09-3.92443835e-13    2
-2.37591504e+04-2.67152365e+01-3.14633439e+00 7.03122692e-02-5.99948828e-05    3
 2.60021921e-08-4.52522129e-12-2.03193740e+04 3.93595186e+01                   4
C6H4O2                  H   4C   6O   2     G    200.00   3500.00 1340.00      1
 9.02248614e+00 2.96818822e-02-1.55447204e-05 3.92075323e-09-3.86404387e-13    2
-1.85718024e+04-2.25961417e+01-1.26066494e+00 6.03778556e-02-4.99058846e-05    3
 2.10158598e-08-3.57578994e-12-1.58159179e+04 3.00236840e+01                   4
C7H7O2                  C   7H   7O   2     G    300.00   3500.00 1420.00      1
 1.76964624e+01 2.58808958e-02-1.00755993e-05 1.78285132e-09-1.17592477e-13    2
 6.43630911e+03-6.45881471e+01-4.45172572e+00 8.82701582e-02-7.59797497e-05    3
 3.27237670e-08-5.56493679e-12 1.27263945e+04 5.00304723e+01                   4
O2C6H4CH3               C   7H   7O   2     G    300.00   3500.00 1300.00      1
 1.57011694e+01 2.91723896e-02-1.27991927e-05 2.73382155e-09-2.31734775e-13    2
 5.63564260e+03-5.46747931e+01-5.21645096e+00 9.35342985e-02-8.70629336e-05    3
 4.08177913e-08-7.55557510e-12 1.10742239e+04 5.17286697e+01                   4
OC6H4CH2                C   7H   6O   1     G    300.00   3500.00 1390.00      1
 1.45795344e+01 2.32519437e-02-8.58329372e-06 1.38947459e-09-7.81466970e-14    2
-5.01093188e+02-5.31869652e+01-4.82277790e+00 7.90859360e-02-6.88358034e-05    3
 3.02875608e-08-5.27564421e-12 4.89274964e+03 4.68072303e+01                   4
C6H5CH2O                C   7H   7O   1     G    300.00   3500.00 1650.00      1
 1.54569227e+01 2.51288522e-02-9.88344275e-06 1.85206220e-09-1.37473827e-13    2
 6.00712849e+03-5.64457004e+01-4.49397764e+00 7.34946712e-02-5.38523691e-05    3
 1.96172850e-08-2.82917425e-12 1.25909256e+04 4.97967788e+01                   4
BZCOOH                  C   7H   8O   2     G    300.00   3500.00 1550.00      1
 1.78036107e+01 3.06807111e-02-1.34555335e-05 2.81495360e-09-2.31878498e-13    2
-1.15055065e+04-6.47324084e+01-3.42659307e+00 8.54683337e-02-6.64758135e-05    3
 2.56193751e-08-3.91001099e-12-4.92414334e+03 4.69952939e+01                   4
C6H5O2                  H   5C   6O   2     G    200.00   3500.00 1360.00      1
 1.04204177e+01 3.01752774e-02-1.55019219e-05 3.86083586e-09-3.77613119e-13    2
 1.18064810e+04-2.92245570e+01-3.03410399e+00 6.97474001e-02-5.91476455e-05    3
 2.52557984e-08-4.31051064e-12 1.54661109e+04 3.98227924e+01                   4
RBBENZ                  C  14H  13          G    300.00   3500.00 1750.00      1
 5.34298872e+01-2.73976091e-03 1.40930518e-05-5.29858386e-09 5.98002536e-13    2
 9.33192271e+03-2.64139662e+02-8.67312060e+00 1.39209971e-01-1.07578147e-04    3
 4.10523491e-08-6.02355932e-12 3.10679755e+04 7.02252758e+01                   4
STILB                   C  14H  12          G    300.00   3500.00 1470.00      1
 3.31295359e+01 3.16424147e-02-7.88066870e-06 4.81370280e-10 4.43949941e-14    2
 1.37146851e+04-1.52659599e+02-1.11031623e+01 1.52003498e-01-1.30698101e-04    3
 5.61808860e-08-9.42831176e-12 2.67190984e+04 7.77787968e+01                   4
HOC6H4CH2               C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353909e-06-2.12687604e-10 1.25840461e-13    2
-3.38086419e+03-4.22339553e+01-6.42956807e+00 9.31830718e-02-9.41722602e-05    3
 5.12938174e-08-1.10712258e-11 1.12339577e+03 5.49833260e+01                   4
OC6H4CH3                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824814e+01 2.40796407e-02-4.51347940e-06-4.25076353e-10 1.44988491e-13    2
-3.97704754e+03-4.00543784e+01-6.60757191e+00 9.15233043e-02-9.24834754e-05    3
 5.05720228e-08-1.09413374e-11 4.82664712e+02 5.62014117e+01                   4
OOC6H4OH                H   5C   6O   3     G    100.00   3500.00 1570.00      1
 2.76569225e+01 2.91346366e-04 5.46428411e-06-2.09157763e-09 2.40972768e-13    2
-1.39658758e+04-1.18517523e+02-4.81896279e-01 7.19826044e-02-6.30305484e-05    3
 2.69932769e-08-4.39037350e-12-5.13028675e+03 2.99287472e+01                   4
C6H4OH                  C   6H   5O   1     G    300.00   3500.00 1170.00      1
 1.35501563e+01 1.98692226e-02-8.43356667e-06 1.70584597e-09-1.35582641e-13    2
 1.32571078e+04-4.75538960e+01-6.19433347e+00 8.73717517e-02-9.49752706e-05    3
 5.10173582e-08-1.06722306e-11 1.78773184e+04 5.08018126e+01                   4
CYC5H10                 C   5H  10          G    300.00   3500.00 1800.00      1
 1.11296301e+01 2.96496234e-02-1.15919105e-05 2.15298805e-09-1.58472912e-13    2
-1.68167420e+04-4.22488373e+01-7.89803624e+00 7.19333263e-02-4.68283297e-05    3
 1.52035137e-08-1.97104591e-12-9.96678208e+03 6.07328622e+01                   4
RCYC5H9                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.66203792e+00 2.81281840e-02-1.16028931e-05 2.36816034e-09-1.95484558e-13    2
 7.45094250e+03-3.11364282e+01-6.79102382e+00 6.46905434e-02-4.20715259e-05    3
 1.36528392e-08-1.76280106e-12 1.33740447e+04 5.79109742e+01                   4
RCYC5H9O2               H   9C   5O   2     g    300.00   3500.00 1490.00      1
 1.41059001e+01 2.93905835e-02-1.10646094e-05 1.87429644e-09-1.16178129e-13    2
-1.11826225e+04-5.13980703e+01-6.20236748e+00 8.39094225e-02-6.59493467e-05    3
 2.64312259e-08-4.23646830e-12-5.13075876e+03 5.46760334e+01                   4
C5H2                    C   5H   2          G    300.00   3500.00 1260.00      1
 1.08586495e+01 8.25356562e-03-3.15379453e-06 5.51063161e-10-3.71272440e-14    2
 7.89908994e+04-3.35264726e+01 1.78531794e+00 3.70577929e-02-3.74445412e-05    3
 1.86943154e-08-3.63697888e-12 8.12773789e+04 1.23440607e+01                   4
C5H3                    C   5H   3          G    300.00   3500.00 1370.00      1
 1.06729929e+01 9.74586302e-03-3.33881730e-06 5.09387247e-10-2.86889361e-14    2
 6.39774214e+04-2.94129104e+01 3.35962353e+00 3.10987662e-02-2.67179083e-05    3
 1.18860739e-08-2.10472664e-12 6.59812846e+04 8.17219633e+00                   4
CYC5H4                  C   5H   4          G    200.00   3500.00 1310.00      1
 6.52292971e+00 1.75112092e-02-7.24525150e-06 1.36813992e-09-9.77801509e-14    2
 6.01459585e+04-1.09295493e+01-1.67820643e+00 4.25528463e-02-3.59188817e-05    3
 1.59603181e-08-2.88254699e-12 6.22946562e+04 3.08507212e+01                   4
C6H2                    C   6H   2          G    200.00   3500.00  700.00      1
 9.95239961e+00 1.43744770e-02-7.32585546e-06 1.80931772e-09-1.74471745e-13    2
 8.06473020e+04-2.49945457e+01-5.39476453e-01 7.43280545e-02-1.35797807e-04    3
 1.24163557e-07-4.38724145e-11 8.21161647e+04 2.18805021e+01                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194523e+01 1.16137832e-02-4.19264521e-06 6.84693068e-10-4.17887563e-14    2
 8.26280760e+04-3.29876543e+01 4.46601449e+00 3.41999583e-02-2.98587533e-05    3
 1.36473739e-08-2.49684195e-12 8.45957836e+04 5.04018538e+00                   4
LC6H4                   C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447675e+01 6.21306704e-03-9.80963831e-07 8.00594547e-11-2.88320672e-15    2
 5.49568894e+04-6.59208083e+01-1.17305610e+00 6.09713718e-02-6.13761529e-05    3
 2.96855443e-08-5.44506792e-12 6.00209374e+04 2.96241244e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076076e+01 1.68261951e-02-6.51181367e-06 1.21158890e-09-8.99428205e-14    2
 5.89425072e+04-3.55373249e+01 1.67614161e-01 5.94226633e-02-6.25597981e-05    3
 3.39881880e-08-7.27779349e-12 6.17104257e+04 2.46218080e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863876e+01 1.90072460e-02-7.30992555e-06 1.31482494e-09-9.21385778e-14    2
 3.55364843e+04-4.09021933e+01-1.05889384e+00 6.36321466e-02-6.08598063e-05    3
 2.98747613e-08-5.80412586e-12 3.90228046e+04 2.94875281e+01                   4
C7H6                    C   7H   6          G    300.00   3500.00 1290.00      1
 1.11282362e+01 2.73165807e-02-1.25329645e-05 2.76951413e-09-2.40721375e-13    2
 3.69620905e+04-3.50553513e+01-3.97785296e+00 7.41571673e-02-6.69987629e-05    3
 3.09172135e-08-5.69570188e-12 4.08594615e+04 4.16694449e+01                   4
C7H5                    C   7H   5          G    300.00   3500.00 1250.00      1
 1.21079560e+01 2.22665290e-02-9.87308079e-06 2.11666746e-09-1.79360812e-13    2
 5.15977924e+04-3.78517160e+01-2.81419579e+00 7.00174146e-02-6.71741435e-05    3
 3.26772342e-08-6.29147417e-12 5.53283304e+04 3.74688223e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155282e-02-1.38949870e-05 2.56768165e-09-1.71519558e-13    2
-2.17187243e+04-3.95715125e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733026e-12-1.73470426e+04 4.54334870e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799877e-06 4.38368234e-10 8.64078966e-14    2
-1.87828963e+04-3.81332334e+01-6.02884975e+00 7.77532977e-02-6.10481841e-05    3
 2.48568442e-08-4.12367417e-12-1.33857950e+04 5.85676633e+01                   4
C6H5C2H                 C   8H   6          G    200.00   3500.00 1280.00      1
 1.52608076e+01 2.33328927e-02-9.12947230e-06 1.67060897e-09-1.19620450e-13    2
 3.14643486e+04-5.61979008e+01-2.98097334e+00 8.03384582e-02-7.59328693e-05    3
 3.64640449e-08-6.91521341e-12 3.61342445e+04 3.63113150e+01                   4
C6H5C2H3                C   8H   8          G    200.00   3500.00 1620.00      1
 2.08689853e+01 1.76153525e-02-4.02709967e-06 7.62333198e-11 4.96213073e-14    2
 7.92336685e+03-8.97908225e+01-4.75261288e+00 8.08785579e-02-6.26041417e-05    3
 2.41820119e-08-3.67040626e-12 1.62247647e+04 4.61791070e+01                   4
C6H5C2H5                C   8H  10          G    200.00   3500.00 1660.00      1
 2.15526224e+01 2.25377527e-02-5.71678491e-06 3.25228910e-10 3.67333515e-14    2
-7.08672427e+03-9.37205827e+01-4.75947977e+00 8.59404087e-02-6.30083415e-05    3
 2.33338862e-08-3.42842587e-12 1.64889367e+03 4.65555372e+01                   4
C6H5C2H2                C   8H   7          G    200.00   3500.00 1520.00      1
 1.92541493e+01 1.80154928e-02-5.00513523e-06 4.35360010e-10 9.55509220e-15    2
 3.83998804e+04-7.81182474e+01-4.29898225e+00 7.99974179e-02-6.61715087e-05    3
 2.72627168e-08-4.40283911e-12 4.55600324e+04 4.53739369e+01                   4
C6H5CHCH3               C   8H   9          G    200.00   3500.00 1700.00      1
 2.17404159e+01 1.87953891e-02-4.10981050e-06 2.63149780e-14 6.24669644e-14    2
 1.18126541e+04-9.21825395e+01-3.04486857e+00 7.71137055e-02-5.55671485e-05    3
 2.01793745e-08-2.90508425e-12 2.02396509e+04 4.05439030e+01                   4
C6H5C2H4                C   8H   9          G    200.00   3500.00 1530.00      1
 1.90733241e+01 2.32393227e-02-7.04814668e-06 8.06136144e-10-1.68209988e-14    2
 1.95612163e+04-7.66267161e+01-3.58296948e+00 8.24714629e-02-6.51188723e-05    3
 2.61092846e-08-4.15132238e-12 2.64940422e+04 4.23117947e+01                   4
C6H4C2H3                C   8H   7          G    200.00   3500.00 1580.00      1
 1.99256075e+01 1.67315530e-02-4.18312961e-06 2.15370099e-10 3.07179808e-14    2
 3.89930312e+04-8.19571079e+01-3.96125911e+00 7.72046330e-02-6.15942816e-05    3
 2.44394849e-08-3.80221157e-12 4.65412811e+04 4.42096620e+01                   4
C6H4C2H                 C   8H   5          G    200.00   3500.00 1410.00      1
 1.60102852e+01 1.80276839e-02-6.10631287e-06 8.89485624e-10-4.39310921e-14    2
 6.01004863e+04-5.91795508e+01-2.59308039e+00 7.08031891e-02-6.22504674e-05    3
 2.74351852e-08-4.75061541e-12 6.53466354e+04 3.69628594e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874483e-03-2.93037073e-06 2.89537319e-10 2.52408504e-16    2
 1.07885460e+05-5.89733616e+01 1.87361690e-01 7.06952486e-02-8.88216497e-05    3
 5.43092096e-08-1.27402363e-11 1.11295389e+05 1.95626384e+01                   4
XYLENE                  C   8H  10          G    200.00   3500.00 1800.00      1
 2.00142025e+01 2.37296570e-02-6.76483884e-06 7.09529215e-10-1.05911395e-14    2
-8.30085767e+03-8.55893311e+01-3.92128796e+00 7.69196357e-02-5.10898211e-05    3
 1.71261893e-08-2.29068282e-12 3.15918887e+02 4.39545364e+01                   4
RXYLENE                 C   8H   9          G    200.00   3500.00 1620.00      1
 2.04972497e+01 2.14206934e-02-5.61362086e-06 3.90126528e-10 2.53125355e-14    2
 1.19614465e+04-8.71674754e+01-3.85447699e+00 8.15484138e-02-6.12874360e-05    3
 2.33011616e-08-3.51034102e-12 1.98514059e+04 4.20634392e+01                   4
INDENE                  C   9H   8          G    200.00   3500.00 1610.00      1
 2.31048443e+01 1.91297591e-02-4.53548120e-06 1.22196710e-10 5.15078704e-14    2
 8.53092089e+03-1.04304478e+02-6.87762290e+00 9.36203608e-02-7.39366630e-05    3
 2.88597461e-08-4.41084452e-12 1.81852753e+04 5.46222708e+01                   4
INDENYL                 H   7C   9          G    300.00   3500.00 1330.00      1
 1.46486993e+01 3.26952593e-02-1.44758057e-05 2.99681991e-09-2.36971392e-13    2
 2.63470874e+04-5.64282180e+01-8.19731515e+00 1.01405077e-01-9.19680816e-05    3
 4.18400660e-08-7.53833343e-12 3.24241273e+04 6.03057978e+01                   4
C10H7                   C  10H   7          G    200.00   3500.00 1490.00      1
 2.12397127e+01 2.27484190e-02-6.96640086e-06 8.04033892e-10-1.68765826e-14    2
 3.76445830e+04-9.11799918e+01-6.45168838e+00 9.70877508e-02-8.18046543e-05    3
 3.42887110e-08-5.63511100e-12 4.58966205e+04 5.34576808e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H7O                  C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C10H6CH3                C  11H   9          G    200.00   3500.00 1530.00      1
 2.52493034e+01 2.50352394e-02-6.91797177e-06 5.80757389e-10 1.70685086e-14    2
 3.22365770e+04-1.13732286e+02-6.94188403e+00 1.09195207e-01-8.94277435e-05    3
 3.65327276e-08-5.85743643e-12 4.20870803e+04 5.52614582e+01                   4
C10H7CH2                C  11H   9          G    200.00   3500.00 1480.00      1
 2.49658354e+01 2.73321443e-02-8.56500981e-06 1.05181516e-09-3.08784850e-14    2
 2.10853669e+04-1.11434350e+02-7.41870774e+00 1.14857936e-01-9.72735830e-05    3
 4.10106319e-08-6.78067861e-12 3.06711917e+04 5.74984546e+01                   4
C10H7CHO                C  11H   8O   1     G    200.00   3500.00 1700.00      1
 3.52801173e+01 1.31180999e-02-5.97608673e-07-9.89256296e-10 1.64132767e-13    2
-1.29136404e+04-1.70276910e+02-6.53399067e+00 1.11504236e-01-8.74089056e-05    3
 3.30543895e-08-4.84228574e-12 1.30315629e+03 5.36397371e+01                   4
C10H7CH3                C  11H  10          G    200.00   3500.00 1700.00      1
 3.19556671e+01 1.89589747e-02-2.92887930e-06-5.41537998e-10 1.30075116e-13    2
-1.51641167e+03-1.52538802e+02-7.17710534e+00 1.11036086e-01-8.41733896e-05    3
 3.13190543e-08-4.55530610e-12 1.17887310e+04 5.70191587e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191869e+01 2.86451308e-02-9.80098219e-06 1.51374083e-09-8.72237945e-14    2
-2.13626711e+04-1.32660114e+02-1.76841814e+00 9.72842531e-02-6.70002508e-05    3
 2.26986551e-08-3.02957300e-12-1.02431333e+04 3.45100483e+01                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936624e+01 3.24954978e-02-1.30480618e-05 2.52260906e-09-1.95492396e-13    2
-2.87396993e+03-1.14905139e+02-1.85059487e+00 9.45938472e-02-6.47966864e-05    3
 2.16887663e-08-2.85745868e-12 7.18596268e+03 3.63350107e+01                   4
C12H8                   C  12H   8          G    200.00   3500.00 1570.00      1
 2.77000801e+01 2.26169409e-02-5.57154154e-06 2.34725134e-10 5.00956725e-14    2
 1.79557632e+04-1.32407942e+02-8.95027490e+00 1.15993641e-01-9.47849497e-05    3
 3.81172764e-08-5.98215771e-12 2.94639746e+04 6.09409166e+01                   4
C12H7                   C  12H   7          G    200.00   3500.00 1550.00      1
 2.72643903e+01 2.07706175e-02-5.09002113e-06 1.94274019e-10 4.95146521e-14    2
 5.03500896e+04-1.28964295e+02-8.21375630e+00 1.12327125e-01-9.36930927e-05    3
 3.83031220e-08-6.09707373e-12 6.13483151e+04 5.77457270e+01                   4
BIPHENYL                C  12H  10          G    200.00   3500.00 1620.00      1
 3.03550325e+01 2.42378629e-02-5.78855002e-06 1.73424746e-10 6.27217930e-14    2
 7.33500914e+03-1.42781766e+02-7.48580974e+00 1.17672041e-01-9.23016780e-05    3
 3.57755350e-08-5.43143103e-12 1.95954420e+04 5.80338349e+01                   4
C12H9                   C  12H   9          G    300.00   3500.00 1430.00      1
 2.37129726e+01 3.27032394e-02-1.16108738e-05 1.80515253e-09-1.00356246e-13    2
 4.00500330e+04-1.02303886e+02-9.58279780e+00 1.25838261e-01-1.09304953e-04    3
 4.73501778e-08-8.06277324e-12 4.95726233e+04 7.02380051e+01                   4
FLUORENE                C  13H  10          G    200.00   3500.00 1580.00      1
 3.04981916e+01 2.54134515e-02-6.12250971e-06 2.13473325e-10 6.26029968e-14    2
 6.42406071e+03-1.44876912e+02-9.12299946e+00 1.25720264e-01-1.01350497e-04    3
 4.03940585e-08-6.29508454e-12 1.89443571e+04 6.43961494e+01                   4
C6H5CH2C6H5             C  13H  12          G    200.00   3500.00 1730.00      1
 3.68978946e+01 2.09448951e-02-2.15140891e-06-1.01983321e-09 1.90993351e-13    2
 1.61235408e+03-1.77722051e+02-9.21937242e+00 1.27574414e-01-9.46047492e-05    3
 3.46076582e-08-4.95748807e-12 1.75689285e+04 7.00449656e+01                   4
C14H10                  C  14H  10          G    200.00   3500.00 1550.00      1
 3.33910328e+01 2.79675689e-02-7.16206047e-06 3.83005680e-10 5.29481034e-14    2
 8.53646106e+03-1.60739744e+02-9.79770356e+00 1.39422372e-01-1.15021548e-04    3
 4.67741830e-08-7.42949985e-12 2.19249693e+04 6.65486198e+01                   4
C14H9                   C  14H   9          G    298.15   3500.00 1380.00      1
 2.51054802e+01 4.12375730e-02-1.71094078e-05 3.35330064e-09-2.55891906e-13    2
 4.20489545e+04-1.12231128e+02-1.15966331e+01 1.47620510e-01-1.32743035e-04    3
 5.92149564e-08-1.03757571e-11 5.21787378e+04 7.66564976e+01                   4
C16H10                  C  16H  10          G    200.00   3500.00 1560.00      1
 3.81807346e+01 2.83119223e-02-6.73305412e-06 1.57165249e-10 8.21178664e-14    2
 9.09208909e+03-1.88517714e+02-1.17161985e+01 1.56252776e-01-1.29753106e-04    3
 5.27298370e-08-8.34298979e-12 2.46599322e+04 7.43946040e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933978e+01 6.96117135e-02-3.71054120e-05 9.43826012e-09-9.32515878e-13    2
 4.61008358e+04-6.54256239e+01-1.33382684e+01 1.64875153e-01-1.52343444e-04    3
 7.13941910e-08-1.34236310e-11 5.34246890e+04 8.34001921e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1170.00      1
 6.79293353e+00 9.36089894e-02-5.25184355e-05 1.38852184e-08-1.40951794e-12    2
 1.04787082e+04-8.65156283e+00-1.16088786e+01 1.56521168e-01-1.33175074e-04    3
 5.98434171e-08-1.12296459e-11 1.47847322e+04 8.30156968e+01                   4
C18H10                  C  18H  10          G    300.00   3500.00 1430.00      1
 3.55205899e+01 2.97059393e-02-5.18578691e-06-7.74972602e-10 2.05763862e-13    2
 1.13998056e+04-1.72584615e+02-1.43149505e+01 1.69106052e-01-1.51409682e-04    3
 6.73946752e-08-1.17120067e-11 2.56527701e+04 8.56679583e+01                   4
C18H9                   C  18H   9          G    300.00   3500.00 1110.00      1
 1.00826780e+01 9.26185738e-02-5.34378516e-05 1.44603235e-08-1.49786389e-12    2
 4.90427510e+04-3.41228885e+01-1.54340436e+01 1.84570724e-01-1.77697514e-04    3
 8.90907512e-08-1.83065188e-11 5.47074632e+04 9.16434687e+01                   4
-9.82259725e+02-1.87789164e+02-1.59101514e+01 1.94323596e-01-1.71453697e-04    3
 7.50992355e-08-1.28697737e-11 1.43320109e+04 8.96934466e+01                   4
-3.16800426e+03-2.10125738e+02-1.45702439e+01 2.15386833e-01-1.89111746e-04    3
 8.32251462e-08-1.44012185e-11 1.27337618e+04 8.12945187e+01                   4
C18H14                  H  14C  18          G    100.00   3500.00  700.00      1
-8.78909816e+00 1.54177573e-01-9.84392858e-05 2.89551422e-08-3.12416385e-12    2
 3.49494076e+04 6.52592557e+01-7.00582263e+00 1.43987427e-01-7.66032589e-05    3
 8.15892605e-09 4.30305619e-12 3.46997490e+04 5.72920318e+01                   4
FC10H10                 H  10C  10          G    290.00   3500.00 1470.00      1
 5.90673294e+00 7.17465912e-02-4.74529572e-05 1.57883693e-08-2.08558667e-12    2
 2.96385223e+04-1.06222118e+01-7.49771949e+00 1.08221292e-01-8.46720393e-05    3
 3.26677716e-08-4.95623333e-12 3.35794313e+04 5.92107542e+01                   4
FC10H10O                H  10C  10O   1     G    290.00   3500.00 1470.00      1
 5.90673294e+00 7.17465912e-02-4.74529572e-05 1.57883693e-08-2.08558667e-12    2
 2.96385223e+04-1.06222118e+01-7.49771949e+00 1.08221292e-01-8.46720393e-05    3
 3.26677716e-08-4.95623333e-12 3.35794313e+04 5.92107542e+01                   4
C9H9                    H   9C   9          G    300.00   3500.00 1420.00      1
 1.65762703e+01 3.32325777e-02-1.27882013e-05 2.22930897e-09-1.43928988e-13    2
 1.59391591e+04-6.61765066e+01-8.97125560e+00 1.05197439e-01-8.88074212e-05    3
 3.79190836e-08-6.42734001e-12 2.31946564e+04 6.60339533e+01                   4
C10H7CH2OOH             C  11H  10O   2     G    200.00   3500.00 1000.00      1
 9.59357183e+00 7.25131639e-02-4.02299427e-05 1.04419273e-08-1.03126748e-12    2
-1.67373561e+03-1.93308213e+01-1.20905039e+01 1.59249467e-01-1.70334397e-04    3
 9.71782303e-08-2.27153432e-11 2.66307954e+03 8.52823095e+01                   4
C10H7CH2O               C  11H   9O   1     G    200.00   3500.00 1000.00      1
 6.19208080e+00 6.85969290e-02-3.75702682e-05 9.69726057e-09-9.55827930e-13    2
 1.63598795e+04-4.97891969e+00-1.25750276e+01 1.43665363e-01-1.50172919e-04    3
 8.47656943e-08-1.97229364e-11 2.01133012e+04 8.55615301e+01                   4
C10H7CH2O2              C  11H   9O   2     G    200.00   3500.00 1000.00      1
 1.10033966e+01 6.55567626e-02-3.57758599e-05 9.18803877e-09-9.01110305e-13    2
 1.54881792e+04-2.80172430e+01-1.29736641e+01 1.61465005e-01-1.79638224e-04    3
 1.05096281e-07-2.48781709e-11 2.02835913e+04 8.76582145e+01                   4
C10H6OH                 C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C10H7C2H5               C  12H  12          G    200.00   3500.00 1710.00      1
 3.70350087e+01 2.11184677e-02-3.34094971e-06-5.61807694e-10 1.38570220e-13    2
-6.26106969e+03-1.80812625e+02-7.78112673e+00 1.25951533e-01-9.52997789e-05    3
 3.52895877e-08-5.10286186e-12 9.06604862e+03 5.94428812e+01                   4
C10H7C2H4               C  12H  11          G    200.00   3500.00 1460.00      1
 2.73240140e+01 3.27963362e-02-1.07965703e-05 1.48242708e-09-6.38934928e-14    2
 2.25065025e+04-1.21828029e+02-6.82202070e+00 1.26347116e-01-1.06910385e-04    3
 4.53700139e-08-7.57889123e-12 3.24771447e+04 5.58289540e+01                   4
C10H7CHCH3              C  12H  11          G    200.00   3500.00 1480.00      1
 2.75888897e+01 3.23001039e-02-1.04831520e-05 1.38976413e-09-5.40501209e-14    2
 1.36246775e+04-1.22421104e+02-6.68326595e+00 1.24927552e-01-1.04362322e-04    3
 4.36776785e-08-7.19727890e-12 2.37692356e+04 5.63583628e+01                   4
C10H6O2                 C  10H   6O   2     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
OC10H6CH2               C  11H   8O   1     G    200.00   3500.00 1000.00      1
 6.19208080e+00 6.85969290e-02-3.75702682e-05 9.69726057e-09-9.55827930e-13    2
 1.63598795e+04-4.97891969e+00-1.25750276e+01 1.43665363e-01-1.50172919e-04    3
 8.47656943e-08-1.97229364e-11 2.01133012e+04 8.55615301e+01                   4
HOC10H6CH2              C  11H   9O   1     G    200.00   3500.00 1000.00      1
 6.19208080e+00 6.85969290e-02-3.75702682e-05 9.69726057e-09-9.55827930e-13    2
 1.63598795e+04-4.97891969e+00-1.25750276e+01 1.43665363e-01-1.50172919e-04    3
 8.47656943e-08-1.97229364e-11 2.01133012e+04 8.55615301e+01                   4
O2C10H6CH3              C  11H   9O   2     G    200.00   3500.00 1000.00      1
 1.10033966e+01 6.55567626e-02-3.57758599e-05 9.18803877e-09-9.01110305e-13    2
 1.54881792e+04-2.80172430e+01-1.29736641e+01 1.61465005e-01-1.79638224e-04    3
 1.05096281e-07-2.48781709e-11 2.02835913e+04 8.76582145e+01                   4
C10H7O2                 C  10H   7O   2     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C9H7O                   C   9H   7O   1     G    300.00   3500.00 1050.00      1
 5.95943049e+00 5.43389701e-02-3.24056700e-05 9.18611701e-09-1.00131985e-12    2
 4.10196259e+03-7.81774446e+00-8.04376203e+00 1.07684465e-01-1.08613520e-04    3
 5.75720538e-08-1.25217810e-11 7.04263302e+03 6.04227829e+01                   4
C9H7OH                  C   9H   8O   1     G    300.00   3500.00 1050.00      1
 5.95943049e+00 5.43389701e-02-3.24056700e-05 9.18611701e-09-1.00131985e-12    2
 4.10196259e+03-7.81774446e+00-8.04376203e+00 1.07684465e-01-1.08613520e-04    3
 5.75720538e-08-1.25217810e-11 7.04263302e+03 6.04227829e+01                   4
C9H6O                   C   9H   6O   1     G    300.00   3500.00 1050.00      1
 5.95943049e+00 5.43389701e-02-3.24056700e-05 9.18611701e-09-1.00131985e-12    2
 4.10196259e+03-7.81774446e+00-8.04376203e+00 1.07684465e-01-1.08613520e-04    3
 5.75720538e-08-1.25217810e-11 7.04263302e+03 6.04227829e+01                   4
C9H6OH                  C   9H   7O   1     G    300.00   3500.00 1050.00      1
 5.95943049e+00 5.43389701e-02-3.24056700e-05 9.18611701e-09-1.00131985e-12    2
 4.10196259e+03-7.81774446e+00-8.04376203e+00 1.07684465e-01-1.08613520e-04    3
 5.75720538e-08-1.25217810e-11 7.04263302e+03 6.04227829e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339062e+01 3.85260822e-02-1.58310821e-05 3.15191459e-09-2.53163787e-13    2
-5.89957979e+03-7.33836419e+01-9.95790328e+00 9.91745477e-02-6.63714701e-05    3
 2.18705768e-08-2.85297798e-12 3.92547162e+03 7.43253244e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194568e+01 4.36180644e-02-1.87773363e-05 3.92059022e-09-3.26702984e-13    2
-2.91866300e+04-7.40611877e+01-1.01006358e+01 1.03218270e-01-6.84441744e-05    3
 2.23157154e-08-2.88158149e-12-1.95313967e+04 7.10947481e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576861e+01 4.50315825e-02-1.97554195e-05 4.21197817e-09-3.57314917e-13    2
-1.09025839e+04-5.35378398e+01-2.75522789e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963371e+01 3.80090295e-02-1.52789389e-05 2.95630099e-09-2.27699217e-13    2
-8.96605283e+03-7.62711275e+01-5.58650157e+00 9.92161261e-02-7.26605920e-05    3
 2.68653231e-08-3.96348393e-12-1.13154446e+03 5.33514397e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777671e+01 3.52558916e-02-1.42493230e-05 2.76058348e-09-2.13045169e-13    2
 6.10938819e+03-7.94713741e+01-1.83523003e+00 8.26181075e-02-5.37178363e-05    3
 1.73785513e-08-2.24331848e-12 1.37820672e+04 3.58790126e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525256e+01 3.24730728e-02-1.15459374e-05 1.79679053e-09-9.97833648e-14    2
-5.30753652e+03-1.13355893e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932248e-08-9.37220079e-12 5.02765510e+03 7.60497478e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623566e-02-8.52218596e-06 1.36123709e-09-7.97159879e-14    2
-5.90596973e+03-6.59480382e+01-8.70136948e+00 9.66875824e-02-8.77887357e-05    3
 3.96542563e-08-7.01685715e-12 1.03797027e+03 6.35339364e+01                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109941e+01 4.74108396e-02-1.82963852e-05 3.42084161e-09-2.57817125e-13    2
-2.68355230e+04-1.31410203e+02-1.02710769e+01 1.32926553e-01-8.95594797e-05    3
 2.98145803e-08-3.92361417e-12-1.29819774e+04 7.68627930e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748171e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565536e-05 2.20632463e-09-1.51941206e-13    2
-9.85314330e+03-1.11161769e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748172e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835938e-02-9.17249483e-06 1.42952537e-09-8.46466190e-14    2
 3.95646505e+03-1.44540610e+02-1.09331574e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619031e+01-7.89283130e-03 1.09697206e-05-3.89489829e-09 4.38586293e-13    2
-1.76924159e+04-2.71823424e+02-1.36343924e+01 1.41210048e-01-1.13282678e-04    3
 4.21245088e-08-5.95299802e-12 6.46225047e+03 9.13157248e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278060e+00 9.04971362e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620333e+01 4.11366392e-02-1.36024110e-05 2.01592783e-09-1.09376626e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278060e+00 9.04971362e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878918e+01 5.29920990e-02-1.98404553e-05 3.55616370e-09-2.54281184e-13    2
-4.56232379e+04-1.22752047e+02-2.17870143e+00 1.22917862e-01-7.81119243e-05    3
 2.51381892e-08-3.25178473e-12-3.42952643e+04 4.75517200e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212692e+01 5.52219738e-02-2.21266526e-05 4.33498891e-09-3.42316503e-13    2
-2.10175171e+04-1.03192977e+02-1.81057271e+00 1.17737178e-01-7.42226562e-05    3
 2.36298050e-08-3.02215208e-12-1.08900540e+04 4.90624204e+01                   4
C10H10                  C  10H  10          G    200.00   3500.00 1650.00      1
 2.68944429e+01 2.21492835e-02-4.82586131e-06-1.98159511e-11 7.73873507e-14    2
 8.93250679e+02-1.25426777e+02-7.42151348e+00 1.05339481e-01-8.04533134e-05    3
 3.05367303e-08-4.55239239e-12 1.22175163e+04 5.73124589e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295230e-05 5.21804510e-09-4.10998519e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710594e-12-1.66984825e+04 5.11161660e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453588e+01 7.53296743e-02-2.79263242e-05 4.92908201e-09-3.44364401e-13    2
-5.61938874e+04-2.43048234e+02-8.95216176e+00 2.21020633e-01-1.60372651e-04    3
 5.84427492e-08-8.45249580e-12-3.63617056e+04 7.69829165e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278371e+01 8.00212238e-02-3.03236334e-05 5.55903617e-09-4.09822554e-13    2
-4.61545210e+04-2.04019480e+02-3.22413374e+00 1.90803381e-01-1.22642098e-04    3
 3.97510601e-08-5.15871477e-12-2.82078115e+04 6.57897857e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414094e+01 6.11045883e-02-2.24641073e-05 3.93182441e-09-2.73349363e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524599e+01 8.54680758e-02-3.36612723e-05 6.38202030e-09-4.82094888e-13    2
-7.78744142e+04-2.24182950e+02-9.93612249e+00 2.29338723e-01-1.69388298e-04    3
 6.32906266e-08-9.42998896e-12-5.96884450e+04 7.82391931e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210237e+01 7.73881688e-02-2.77557896e-05 4.69678103e-09-3.12959243e-13    2
-7.08514663e+04-2.24842855e+02-3.64057977e+00 1.96191732e-01-1.26758759e-04    3
 4.13645475e-08-5.40570458e-12-5.16052891e+04 6.45024954e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971791e+01 4.89478938e-02-1.82737062e-05 3.23575201e-09-2.26811842e-13    2
-3.12534582e+04-1.16784058e+02-2.31417710e+00 1.16973130e-01-7.49614029e-05    3
 2.42311952e-08-3.14284563e-12-2.02333700e+04 4.88909878e+01                   4
IC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414094e+01 6.11045883e-02-2.24641073e-05 3.93182441e-09-2.73349363e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
IC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295230e-05 5.21804510e-09-4.10998519e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710594e-12-1.66984825e+04 5.11161660e+01                   4
C10H16                  C  10H  16          G    300.00   3500.00 1800.00      1
 2.89286921e+01 4.33698641e-02-1.66040771e-05 3.00058011e-09-2.14826944e-13    2
-2.62354027e+04-1.44986840e+02-1.64117649e+01 1.44126435e-01-1.00567886e-04    3
 3.40982872e-08-4.53395293e-12-9.91283823e+03 1.00405171e+02                   4
C10H15                  C  10H  15          G    300.00   3500.00 1770.00      1
 3.20501672e+01 3.53882361e-02-1.22004701e-05 1.87186214e-09-1.05121248e-13    2
-9.38259390e+03-1.63611897e+02-1.67888481e+01 1.45758892e-01-1.05734924e-04    3
 3.71014118e-08-5.08104634e-12 7.90641753e+03 9.98941988e+01                   4
C6H5C4H9                C  10H  14          G    300.00   3500.00 1620.00      1
 2.20508088e+01 4.25105888e-02-1.68597965e-05 3.21476378e-09-2.44036713e-13    2
-1.30455855e+04-9.17623601e+01-5.81141602e+00 1.11306205e-01-8.05594416e-05    3
 2.94286095e-08-4.28938328e-12-4.01822468e+03 5.60982344e+01                   4
RC6H5C4H8               C  10H  13          G    300.00   3500.00 1650.00      1
 2.28150862e+01 3.94891782e-02-1.56943357e-05 2.97948809e-09-2.24328827e-13    2
 4.22313026e+03-9.69374623e+01-3.49464028e+00 1.03270333e-01-7.36772040e-05    3
 2.64069096e-08-3.77393815e-12 1.29053400e+04 4.31670204e+01                   4
C6H5C4H7-3              C  10H  12          G    300.00   3500.00 1480.00      1
 1.62604546e+01 4.74926138e-02-2.11208270e-05 4.52915802e-09-3.83727993e-13    2
 2.53220324e+03-5.97390118e+01-5.26848595e+00 1.05678940e-01-8.00934545e-05    3
 3.10934047e-08-4.87093182e-12 8.90476965e+03 5.25659324e+01                   4
CH2OHCH2OH              C   2H   6O   2     G    300.00   3500.00 1510.00      1
 8.58229286e+00 1.47365725e-02-4.87454255e-06 7.03407966e-10-3.54291380e-14    2
-5.09140292e+04-1.61663169e+01-4.19778978e-01 3.85831204e-02-2.85631663e-05    3
 1.11619615e-08-1.76697774e-12-4.81954035e+04 3.09733167e+01                   4
GLYCEROL                C   3H   8O   3     G    300.00   3500.00 1260.00      1
 1.38765805e+01 2.06689859e-02-7.56631173e-06 1.26540495e-09-8.07916650e-14    2
-7.51651919e+04-3.83652419e+01 3.56065369e+00 5.34179600e-02-4.65531857e-05    3
 2.18933806e-08-4.17364397e-12-7.25655783e+04 1.37872736e+01                   4
C3H4O3                  C   3H   4O   3     G    300.00   3500.00 1710.00      1
 1.37242810e+01 1.08811110e-02-3.70124855e-06 5.78901441e-10-3.43205819e-14    2
-5.77802807e+04-3.99570073e+01 2.17563103e+00 3.78954970e-02-2.73980784e-05    3
 9.81743158e-09-1.38498288e-12-5.38306424e+04 2.19543274e+01                   4
FURFURAL                C   5H   4O   2     G    300.00   3500.00 1430.00      1
 1.05158963e+01 2.23224229e-02-1.09267096e-05 2.56683236e-09-2.34844996e-13    2
-2.33303219e+04-2.94000375e+01-1.81996645e+00 5.68283326e-02-4.71217198e-05    3
 1.94409630e-08-3.18486783e-12-1.98022652e+04 3.45255921e+01                   4
FURAN                   C   4H   4O   1     G    300.00   3500.00 1250.00      1
 8.37486468e+00 1.95634451e-02-9.90167118e-06 2.37694381e-09-2.20517697e-13    2
-9.41817580e+03-2.52053385e+01-7.59507782e+00 7.06672611e-02-7.12262504e-05    3
 3.50833860e-08-6.76180614e-12-5.42569018e+03 5.54039923e+01                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   3500.00 1590.00      1
 1.05858550e+01 1.29956017e-02-4.76361254e-06 7.49449812e-10-3.96847799e-14    2
 3.10513348e+03-2.93262371e+01 1.05972039e+00 3.69607201e-02-2.73722149e-05    3
 1.02289476e-08-1.53017186e-12 6.13444428e+03 2.10494483e+01                   4
C4H3O                   C   4H   3O   1     G    300.00   3500.00 1240.00      1
 8.44125907e+00 1.62911135e-02-8.34126433e-06 2.01436765e-09-1.87394602e-13    2
 1.94535776e+04-2.27855079e+01-5.90872254e+00 6.25813768e-02-6.43375505e-05    3
 3.21198979e-08-6.25705795e-12 2.30123730e+04 4.95317027e+01                   4
MEFU2                   C   5H   6O   1     G    300.00   3500.00 1260.00      1
 5.16398170e+00 3.29529080e-02-1.68209195e-05 4.03716052e-09-3.55511368e-13    2
-1.31841670e+04-2.67616715e+00-3.74149805e+00 6.12242723e-02-5.04773056e-05    3
 2.18447722e-08-3.88876765e-12-1.09399861e+04 4.23457855e+01                   4
DMF-3YL                 C   6H   7O   1     G    300.00   3500.00 1620.00      1
 1.41703395e+01 2.18230092e-02-7.69511406e-06 1.17891300e-09-6.12376633e-14    2
 1.19557792e+04-4.86583490e+01-1.12307985e+00 5.95845385e-02-4.26594930e-05    3
 1.55675463e-08-2.28170577e-12 1.69108471e+04 3.25015044e+01                   4
C6H10O5                 C   6H  10O   5     G    300.00   3500.00 1220.00      1
 1.54889719e+01 4.96354386e-02-2.45944508e-05 5.82332583e-09-5.35665861e-13    2
-1.09180509e+05-4.81819838e+01-7.95116462e+00 1.26488345e-01-1.19085729e-04    3
 5.74579043e-08-1.11165221e-11-1.03461116e+05 6.95642163e+01                   4
C6H8O4                  C   6H   8O   4     G    300.00   3500.00 1300.00      1
 1.58073709e+01 3.77998882e-02-1.77241312e-05 3.97560136e-09-3.49009860e-13    2
-7.78788467e+04-5.15128322e+01-4.55493836e+00 1.00453147e-01-9.00163533e-05    3
 4.10485358e-08-7.47842033e-12-7.25846463e+04 5.20658817e+01                   4
C6H6O3                  C   6H   6O   3     G    300.00   3500.00 1770.00      1
 1.98638073e+01 1.79335016e-02-5.95408858e-06 8.93593938e-10-4.95459879e-14    2
-4.95264845e+04-7.44496694e+01 7.10718581e-01 6.12173180e-02-4.26352889e-05    3
 1.47094886e-08-2.00094354e-12-4.27462910e+04 2.88889342e+01                   4
C5H8O4                  C   5H   8O   4     G    300.00   3500.00 1230.00      1
 1.19601536e+01 3.99450842e-02-1.95947372e-05 4.60940116e-09-4.22302288e-13    2
-8.26385858e+04-2.91875209e+01-6.95683232e+00 1.01463738e-01-9.46174852e-05    3
 4.52721372e-08-8.68708604e-12-7.79850073e+04 6.59920851e+01                   4
CATECHOL                C   6H   6O   2     G    300.00   3500.00 1150.00      1
 1.43499798e+01 2.44086034e-02-1.04210955e-05 2.01938915e-09-1.47232753e-13    2
-3.94515399e+04-4.76262861e+01-5.49815264e+00 9.34455857e-02-1.00469333e-04    3
 5.42212661e-08-1.14954669e-11-3.48864694e+04 5.09034930e+01                   4
GUAIACOL                C   7H   8O   2     G    300.00   3500.00 1000.00      1
 9.99301702e+00 4.50609511e-02-2.36180854e-05 5.74986028e-09-5.33615163e-13    2
-3.55531885e+04-2.30989094e+01-7.52910625e+00 1.15149444e-01-1.28750825e-04    3
 7.58383534e-08-1.80557384e-11-3.20487639e+04 6.14352066e+01                   4
SALICALD                C   7H   6O   2     G    300.00   3500.00 1580.00      1
 2.23242869e+01 1.54051239e-02-2.83991520e-06-4.41655604e-10 1.22876781e-13    2
-3.64536802e+04-8.95534660e+01-5.00623399e+00 8.45963160e-02-6.85277558e-05    3
 2.72747329e-08-4.26262772e-12-2.78172356e+04 5.48021581e+01                   4
VANILLIN                C   8H   8O   3     G    300.00   3500.00 1260.00      1
 1.36544657e+01 4.84143206e-02-2.42641773e-05 5.50487741e-09-4.76001842e-13    2
-5.18855417e+04-3.54575763e+01-4.86637434e+00 1.07210638e-01-9.42597934e-05    3
 4.25395949e-08-7.82416008e-12-4.72182901e+04 5.81751540e+01                   4
C8H6O3                  C   8H   6O   3     G    300.00   3500.00 1000.00      1
 4.59308938e+00 6.23299053e-02-3.47374653e-05 8.74937512e-09-8.39789340e-13    2
-4.48191760e+04 1.51136268e+01-8.47052157e+00 1.14584349e-01-1.13119131e-04    3
 6.10038189e-08-1.39034003e-11-4.22064538e+04 7.81379982e+01                   4
C6H5OCH3                C   7H   8O   1     G    300.00   3500.00 1380.00      1
 1.25085136e+01 3.49906122e-02-1.63096082e-05 3.64836833e-09-3.19988393e-13    2
-1.52038795e+04-4.20406498e+01-5.29461551e+00 8.65938851e-02-7.24001222e-05    3
 3.07452350e-08-5.22884105e-12-1.02902159e+04 4.95832512e+01                   4
C7H6O3                  C   7H   6O   3     G    300.00   3500.00 1000.00      1
 9.61003482e+00 4.63126508e-02-2.49854466e-05 6.23131070e-09-5.96782041e-13    2
-5.28813088e+04-1.46625767e+01-7.07010661e+00 1.13033217e-01-1.25066295e-04    3
 7.29518764e-08-1.72769235e-11-4.95452805e+04 6.58094637e+01                   4
RC7H5O3                 C   7H   5O   3     G    300.00   3500.00 1000.00      1
 1.03519979e+01 4.06949751e-02-2.16398121e-05 5.16863286e-09-4.69580368e-13    2
-3.48541025e+04-1.78724723e+01-6.94106369e+00 1.09867221e-01-1.25398181e-04    3
 7.43408790e-08-1.77626419e-11-3.13954902e+04 6.55565533e+01                   4
C24H28O4                C  24H  28O   4     G    300.00   3500.00 1080.00      1
 1.29252083e+01 8.11297204e-02-4.64957343e-05 1.23575596e-08-1.22239418e-12    2
-7.66058401e+03-2.94388917e+00 3.08710551e+00 1.17567138e-01-9.71032588e-05    3
 4.35967723e-08-8.45369342e-12-5.53555381e+03 4.52764204e+01                   4
RSALICPH                C   7H   5O   2     G    300.00   3500.00 1000.00      1
 6.00653618e+00 4.55336023e-02-2.51852438e-05 6.39158463e-09-6.19568356e-13    2
 4.68000597e+02 2.82366668e+00-8.00629363e+00 1.01584922e-01-1.09262223e-04    3
 6.24429039e-08-1.46323982e-11 3.27056656e+03 7.04274704e+01                   4
RGUAIPH                 C   7H   7O   2     G    300.00   3500.00 1000.00      1
 1.03288605e+01 4.15815436e-02-2.20221230e-05 5.39151185e-09-5.01575209e-13    2
-4.91455279e+03-2.20047760e+01-7.23884832e+00 1.11852379e-01-1.27428376e-04    3
 7.56623473e-08-1.80692841e-11-1.40101102e+03 6.27492641e+01                   4
C6H4OCH3                C   7H   7O   1     G    300.00   3500.00 1000.00      1
 6.14038338e+00 4.52741698e-02-2.46495239e-05 6.30633007e-09-6.15603035e-13    2
 1.78813933e+04-4.35386646e+00-8.02841875e+00 1.01949378e-01-1.09662337e-04    3
 6.29815386e-08-1.47844052e-11 2.07151538e+04 6.40024135e+01                   4
RCATEPH                 C   6H   5O   2     G    300.00   3500.00 1000.00      1
 1.18218909e+01 2.70911128e-02-1.34162451e-05 3.08575096e-09-2.72412002e-13    2
-7.82412457e+03-3.10506064e+01-7.41421160e+00 1.04035523e-01-1.28832860e-04    3
 8.00301608e-08-1.95085145e-11-3.97690408e+03 6.17524685e+01                   4
CYC5H4CO                C   6H   4O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658729e-02-6.67332776e-06 1.12237516e-09-7.10809492e-14    2
 1.54076839e+04-4.72500521e+01-4.80707079e+00 7.32685627e-02-6.95172935e-05    3
 3.28617518e-08-6.08232653e-12 2.02256542e+04 4.58618545e+01                   4
NO                      N   1O   1          G    200.00   3500.00  800.00      1
 2.84621514e+00 2.06354046e-03-1.06904715e-06 2.65706521e-10-2.54948672e-14    2
 1.00671113e+04 8.61842850e+00 4.25026596e+00-4.95671364e-03 1.20939293e-05    3
-1.07034405e-08 3.40236358e-12 9.84246312e+03 2.15799981e+00                   4
N2O                     N   2O   1          G    200.00   3500.00 1420.00      1
 4.85543722e+00 2.58052440e-03-9.33594196e-07 1.54088463e-10-9.24862861e-15    2
 8.05595827e+03-2.39060855e+00 2.51620681e+00 9.16990584e-03-7.89420840e-06    3
 3.42198245e-09-5.84582078e-13 8.72029970e+03 9.71509320e+00                   4
NO2                     N   1O   2          G    200.00   3500.00 1800.00      1
 4.19813794e+00 3.78881378e-03-2.08226003e-06 5.53837970e-10-5.45690377e-14    2
 2.49824368e+03 3.49647574e+00 2.86592221e+00 6.74929318e-03-4.54932620e-06    3
 1.46756618e-09-1.81475734e-13 2.97784134e+03 1.07067052e+01                   4
HNO                     H   1N   1O   1     G    200.00   3500.00  700.00      1
 2.88552845e+00 3.71507602e-03-9.89194574e-07 1.60505676e-10-1.61198692e-14    2
 1.18465422e+04 9.10108585e+00 4.47186928e+00-5.34972868e-03 1.84353869e-05    3
-1.83390957e-08 6.59088064e-12 1.16244545e+04 2.01371640e+00                   4
HNO2                    H   1N   1O   2     G    200.00   3500.00  700.00      1
 1.72007297e+00 1.13464166e-02-6.67663344e-06 1.82835451e-09-1.88889111e-13    2
-6.26025905e+03 1.58192354e+01 3.09881792e+00 3.46787404e-03 1.02059578e-05    3
-1.42503038e-08 5.55348885e-12-6.45328334e+03 9.65935177e+00                   4
HONO                    H   1N   1O   2     G    200.00   3500.00 1450.00      1
 5.99816567e+00 3.29505604e-03-1.07588927e-06 1.49768833e-10-6.76019596e-15    2
-1.16909495e+04-5.24156198e+00 2.71684795e+00 1.23469670e-02-1.04399351e-05    3
 4.45507726e-09-7.49054752e-13-1.07393674e+04 1.18081173e+01                   4
HONO2                   H   1N   1O   3     G    200.00   3500.00 1480.00      1
 8.72243659e+00 3.29016496e-03-9.97289211e-07 9.83685339e-11 7.21002272e-16    2
-1.96262630e+04-2.01737896e+01 1.12599207e+00 2.38210961e-02-2.18056654e-05    3
 9.47151094e-09-1.58258008e-12-1.73777154e+04 1.94527900e+01                   4
N2H2                    N   2H   2          G    200.00   3500.00  700.00      1
 1.61507706e+00 8.37729351e-03-2.70267465e-06 3.47805192e-10-1.28897309e-14    2
 2.32788099e+04 1.47543853e+01 4.76517118e+00-9.62324433e-03 3.58699064e-05    3
-3.63879863e-08 1.31070358e-11 2.28377967e+04 6.80561766e-01                   4
H2NN                    N   2H   2          G    200.00   3500.00  700.00      1
 1.58440836e+00 9.29486030e-03-4.50990677e-06 1.06229464e-09-9.86121900e-14    2
 3.53712259e+04 1.46993890e+01 4.53650991e+00-7.57429138e-03 3.16382754e-05    3
-3.33645455e-08 1.21966879e-11 3.49579317e+04 1.51014616e+00                   4
HNNO                    H   1O   1N   2     G    300.00   3500.00 1360.00      1
 4.88500308e+00 5.60936901e-03-2.60717829e-06 5.93839035e-10-5.41495113e-14    2
 2.58926738e+04 6.01979999e-01 2.29344826e+00 1.32315890e-02-1.10140386e-05    3
 4.71484900e-09-8.11688108e-13 2.65975767e+04 1.39015974e+01                   4
NH2NO                   N   2H   2O   1     G    300.00   3500.00 1800.00      1
 5.77099802e+00 9.34065402e-03-4.91077891e-06 1.15317893e-09-1.04142499e-13    2
 6.27743878e+03-6.42402625e+00 1.47077476e+00 1.88967057e-02-1.28741553e-05    3
 4.10257760e-09-5.13781203e-13 7.82551915e+03 1.68496791e+01                   4
NH2OH                   N   1H   3O   1     G    200.00   3500.00 1140.00      1
 3.89950480e+00 8.10759690e-03-2.78780416e-06 4.26313677e-10-2.40531456e-14    2
-6.86348423e+03 3.69890739e+00 2.36719772e+00 1.34841130e-02-9.86216739e-06    3
 4.56336820e-09-9.31301944e-13-6.51411822e+03 1.12921788e+01                   4
HNOH                    H   2N   1O   1     G    200.00   3500.00 1800.00      1
 3.80328699e+00 5.45108878e-03-2.14629752e-06 4.23543078e-10-3.43983588e-14    2
 1.05861530e+04 4.48881947e+00 2.57438367e+00 8.18198504e-03-4.42204441e-06    3
 1.26641230e-09-1.51463528e-13 1.10285582e+04 1.11399006e+01                   4
NH3                     H   3N   1          G    200.00   3500.00  700.00      1
 2.51781806e+00 5.95384021e-03-2.00551774e-06 3.21049856e-10-1.88806102e-14    2
-6.46278678e+03 7.18902506e+00 4.05091142e+00-2.80669327e-03 1.67670540e-05    3
-1.75575899e-08 6.36634787e-12-6.67741985e+03 3.39551804e-01                   4
N2H4                    N   2H   4          G    200.00   3500.00 1780.00      1
 6.33303156e+00 6.50860837e-03-1.68647513e-06 1.37724242e-10 3.10842629e-15    2
 8.61374481e+03-1.06617323e+01 1.71754283e+00 1.68804931e-02-1.04268275e-05    3
 3.41126444e-09-4.56658456e-13 1.02568588e+04 1.42666853e+01                   4
N                       N   1               G    200.00   3500.00 1800.00      1
 2.42215558e+00 1.52655402e-04-9.87414150e-08 2.32518158e-11-1.22034407e-15    2
 5.61344054e+04 4.62162566e+00 2.50554288e+00-3.26497078e-05 5.56795096e-08    3
-3.39411193e-11 6.72311912e-15 5.61043859e+04 4.17031620e+00                   4
NO3                     N   1O   3          G    200.00   3500.00 1380.00      1
 7.84336636e+00 1.94266904e-03-6.08797820e-07 6.42446445e-11-1.29735613e-16    2
 5.97435425e+03-1.61838197e+01 7.80028063e-01 2.24161134e-02-2.28625417e-05    3
 1.08148455e-08-1.94770236e-12 7.92383562e+03 2.01676893e+01                   4
NH                      N   1H   1          G    200.00   3500.00 1670.00      1
 2.48662839e+00 1.81565444e-03-7.12541166e-07 1.51936873e-10-1.23899449e-14    2
 4.24864648e+04 7.43461547e+00 3.66298286e+00-1.00196106e-03 1.81825120e-06    3
-8.58359483e-10 1.38852024e-13 4.20935624e+04 1.15612276e+00                   4
NNH                     N   2H   1          G    200.00   3500.00  740.00      1
 2.70691639e+00 4.73245691e-03-2.26389292e-06 5.23129547e-10-4.76635006e-14    2
 2.90245412e+04 1.03117271e+01 4.29167562e+00-3.83380923e-03 1.51001601e-05    3
-1.51201614e-08 5.23723210e-12 2.87899969e+04 3.14335891e+00                   4
NH2                     N   1H   2          G    200.00   3500.00 1280.00      1
 2.55273412e+00 3.54675597e-03-1.12718085e-06 1.61534507e-10-6.97197514e-15    2
 2.15912601e+04 8.13032012e+00 4.10678625e+00-1.30965693e-03 4.56392802e-06    3
-2.80258469e-09 5.71957556e-13 2.11934228e+04 2.49283504e-01                   4
H2NO                    N   1H   2O   1     G    200.00   3500.00  700.00      1
 2.72801504e+00 7.40936630e-03-3.46220929e-06 8.08344164e-10-7.54853118e-14    2
 6.86495538e+03 9.84388852e+00 3.66110547e+00 2.07742097e-03 7.96338783e-06    3
-1.00731769e-08 3.81077221e-12 6.73432272e+03 5.67507654e+00                   4
N2H3                    N   2H   3          G    200.00   3500.00 1800.00      1
 4.54460800e+00 6.62772042e-03-2.15038229e-06 3.20318188e-10-1.81983291e-14    2
 2.50493358e+04-4.68168818e-02 2.12003669e+00 1.20156567e-02-6.64032916e-06    3
 1.98326147e-09-2.49162674e-13 2.59221815e+04 1.30754688e+01                   4
HCN                     H   1C   1N   1     G    200.00   3500.00  780.00      1
 3.49786301e+00 3.76915270e-03-1.51027204e-06 3.01080816e-10-2.43629369e-14    2
 1.43955802e+04 3.23683734e+00 2.24572677e+00 1.01903642e-02-1.38587556e-05    3
 1.08553403e-08-3.40713841e-12 1.45909135e+04 8.96656341e+00                   4
HNC                     H   1N   1C   1     G    200.00   3500.00  700.00      1
 4.41179651e+00 2.12707775e-03-4.71968008e-07 1.02354109e-12 7.69770096e-15    2
 2.16589078e+04-1.07356913e+00 2.73172542e+00 1.17274840e-02-2.10442671e-05    3
 1.95936894e-08-6.98968295e-12 2.18941178e+04 6.43256347e+00                   4
HNCO                    H   1N   1C   1O   1G    200.00   3500.00 1050.00      1
 4.68274059e+00 5.27517046e-03-2.30255409e-06 4.91740802e-10-4.20405691e-14    2
-1.59709573e+04 2.61731788e-01 2.23902625e+00 1.45845584e-02-1.56016797e-05    3
 8.93563010e-09-2.05249040e-12-1.54577773e+04 1.21704701e+01                   4
HCNO                    H   1N   1C   1O   1G    200.00   3500.00  780.00      1
 4.79767988e+00 6.41431463e-03-3.21741496e-06 7.84733932e-10-7.49876223e-14    2
 1.84217969e+04-2.20789645e+00 6.69823293e-01 2.75828100e-02-4.39260598e-05    3
 3.55784475e-08-1.12268189e-11 1.90657425e+04 1.66810126e+01                   4
HOCN                    H   1N   1C   1O   1G    200.00   3500.00 1260.00      1
 5.08605507e+00 4.40745638e-03-1.67135017e-06 3.00184383e-10-2.12769828e-14    2
-3.69516510e+03-1.53122287e+00 2.95277827e+00 1.11797637e-02-9.73362079e-06    3
 4.56593603e-09-8.67656279e-13-3.15757934e+03 9.25362984e+00                   4
CH2NO                   C   1H   2N   1O   1G    200.00   3500.00 1800.00      1
 3.20402663e+00-6.01464842e-03 5.38459530e-05-6.82208893e-08 2.71923018e-11    2
 2.61694738e+04 1.15885396e+01 8.41613784e+00-1.75971178e-02 6.34980108e-05    3
-7.17957255e-08 2.76888068e-11 2.42931138e+04-1.66204936e+01                   4
CH3NO                   C   1H   3N   1O   1G    200.00   3500.00  700.00      1
 1.71612018e+00 1.65151446e-02-8.81735210e-06 2.26713780e-09-2.25490383e-13    2
 7.35980364e+03 1.71612004e+01 4.07025676e+00 3.06293560e-03 2.00088101e-05    3
-2.51863500e-08 9.57932670e-12 7.03022452e+03 6.64351378e+00                   4
CH3NO2                  C   1H   3N   1O   2G    200.00   3500.00 1800.00      1
 5.69934620e+00 1.38065607e-02-6.43453311e-06 1.45264682e-09-1.30225206e-13    2
-1.27635731e+04-5.01015009e+00 5.58676790e-01 2.52302705e-02-1.59542913e-05    3
 4.97848318e-09-6.19924700e-13-1.09129321e+04 2.28122252e+01                   4
CH3ONO                  C   1H   3O   2N   1G    200.00   3500.00  700.00      1
 2.81666881e+00 1.89749543e-02-1.04049679e-05 2.71704314e-09-2.72624829e-13    2
-9.44747973e+03 1.52094758e+01 5.07409808e+00 6.07535848e-03 1.72370231e-05    3
-2.36086626e-08 9.12941293e-12-9.76351983e+03 5.12385293e+00                   4
CH3ONO2                 C   1H   3N   1O   3G    200.00   3500.00 1800.00      1
 1.20582369e+01 7.66565557e-03-2.49975436e-06 3.22039324e-10-1.19527488e-14    2
-2.00738863e+04-3.71551340e+01 2.05585055e+00 2.98931809e-02-2.10226921e-05    3
 7.18238664e-09-9.64778764e-13-1.64730272e+04 1.69798677e+01                   4
CH3CN                   C   2H   3N   1     G    200.00   3500.00  700.00      1
 2.04918664e+00 1.63166629e-02-8.45703420e-06 2.11771927e-09-2.06450509e-13    2
 7.64801686e+03 1.30927474e+01 3.05185721e+00 1.05871167e-02 3.82056461e-06    3
-9.57523198e-09 3.96960351e-12 7.50764298e+03 8.61306899e+00                   4
CN                      C   1N   1          G    200.00   3500.00  890.00      1
 2.80498942e+00 1.99013249e-03-1.04863794e-06 2.95566162e-10-3.14165336e-14    2
 5.18669927e+04 7.89927658e+00 3.76469138e+00-2.32313475e-03 6.22091360e-06    3
-5.14979080e-09 1.49817812e-12 5.16961658e+04 3.38110710e+00                   4
NCN                     C   1N   2          G    200.00   3500.00 1540.00      1
 6.26178527e+00 8.14604744e-04-6.32168058e-08-5.68978567e-11 1.02757866e-14    2
 5.13388447e+04-9.55046103e+00 2.82367216e+00 9.74476868e-03-8.76142843e-06    3
 3.70856172e-09-6.01000119e-13 5.23977836e+04 8.52096412e+00                   4
NCO                     N   1C   1O   1     G    200.00   3500.00 1630.00      1
 5.49723499e+00 1.70371834e-03-5.14809903e-07 5.30240357e-11-1.05670805e-16    2
 1.33777864e+04-4.53940223e+00 2.90100726e+00 8.07482934e-03-6.37779548e-06    3
 2.45097315e-09-3.67889277e-13 1.42241566e+04 9.25436079e+00                   4
HNCN                    C   1H   1N   2     G    200.00   3500.00 1460.00      1
 5.71563435e+00 3.59039536e-03-1.19666899e-06 1.72409983e-10-8.44530525e-15    2
 3.58827351e+04-4.39973155e+00 3.04255635e+00 1.09138967e-02-8.72081421e-06    3
 3.60809273e-09-5.96747146e-13 3.66632738e+04 9.50791468e+00                   4
H2CN                    C   1H   2N   1     G    200.00   3500.00  700.00      1
 2.09516104e+00 9.19258718e-03-4.75958105e-06 1.19375090e-09-1.16674695e-13    2
 2.77113212e+04 1.25272169e+01 3.31830755e+00 2.20317854e-03 1.02177232e-05    3
-1.30703484e-08 4.97764647e-12 2.75400807e+04 7.06250774e+00                   4
HCNH                    C   1H   2N   1     G    200.00   3500.00  700.00      1
 2.20517225e+00 9.23158578e-03-4.92876098e-06 1.27407702e-09-1.27539972e-13    2
 3.17668288e+04 1.24496856e+01 2.93126392e+00 5.08249047e-03 3.96215754e-06    3
-7.19346443e-09 2.89658197e-12 3.16651760e+04 9.20569165e+00                   4
C2N2                    C   2N   2          G    200.00   3500.00  700.00      1
 5.66789416e+00 5.81681879e-03-2.89262850e-06 6.98368847e-10-6.54524517e-14    2
 3.52445641e+04-4.84945633e+00 2.74684249e+00 2.25085426e-02-3.86606081e-05    3
 3.47631114e-08-1.22314319e-11 3.56535113e+04 8.20106351e+00                   4
CH2CN                   C   2H   2N   1     G    300.00   3500.00 1350.00      1
 4.88864306e+00 8.97936886e-03-4.42991056e-06 1.04146331e-09-8.86722374e-14    2
 2.97135249e+04-5.23788565e-01 3.14472180e+00 1.41465430e-02-1.01712151e-05    3
 3.87667544e-09-6.13711521e-13 3.01843836e+04 8.41298223e+00                   4
CH2NH                   C   1H   3N   1     G    200.00   3500.00  700.00      1
 5.80669265e-01 1.46544725e-02-7.73860026e-06 1.97648489e-09-1.95880938e-13    2
 9.93682812e+03 1.93649676e+01 3.61447523e+00-2.68156156e-03 2.94100442e-05    3
-3.34031765e-08 1.24397124e-11 9.51209529e+03 5.81069013e+00                   4
CH3NH2                  C   1H   5N   1     G    200.00   3500.00  700.00      1
 1.20284786e-02 2.20167260e-02-1.17795638e-05 3.04373591e-09-3.04205303e-13    2
-3.36839831e+03 2.22359932e+01 3.27259122e+00 3.38493895e-03 2.81456942e-05    3
-3.49803194e-08 1.32758144e-11-3.82487709e+03 7.66862375e+00                   4
CH2NH2                  C   1H   4N   1     G    200.00   3500.00 1610.00      1
 5.12514693e+00 8.47270266e-03-2.64074178e-06 3.52691280e-10-1.53029317e-14    2
 1.56058530e+04-3.27656794e+00 1.70381408e+00 1.69729085e-02-1.05601882e-05    3
 3.63196517e-09-5.24506951e-13 1.67075222e+04 1.48587410e+01                   4
CH3NH                   C   1H   4N   1     G    200.00   3500.00  700.00      1
 1.06266679e+00 1.68343860e-02-8.55523919e-06 2.12514555e-09-2.06816968e-13    2
 2.05050909e+04 1.75854917e+01 3.52441786e+00 2.76723702e-03 2.15886516e-05    3
-2.65833218e-08 1.00462071e-11 2.01604458e+04 6.58701073e+00                   4
DMF                     C   6H   8O   1     G    300.00   3500.00 1590.00      1
 1.38889506e+01 2.49736923e-02-8.98421019e-06 1.42738237e-09-7.97717940e-14    2
-2.20872034e+04-4.94041110e+01-2.31533181e+00 6.57391826e-02-4.74422199e-05    3
 1.75523340e-08-2.61514155e-12-1.69342416e+04 3.62866615e+01                   4
CH3OCH3                 C   2H   6O   1     G    300.00   3500.00 1800.00      1
 4.75054344e+00 1.85969149e-02-7.67398366e-06 1.52676542e-09-1.21721364e-13    2
-2.48946055e+04-1.32909286e+00 8.26271488e-01 2.73175193e-02-1.49411539e-05    3
 4.21830997e-09-4.95546995e-13-2.34818676e+04 1.99098856e+01                   4
CH3OCH2                 C   2H   5O   1     G    300.00   3500.00 1800.00      1
 4.38698061e+00 1.62462172e-02-6.72869594e-06 1.35709490e-09-1.09478907e-13    2
-2.38681592e+03 3.59290257e+00 1.56125470e+00 2.25256081e-02-1.19615217e-05    3
 3.29517851e-09-3.78657186e-13-1.36955459e+03 1.88863207e+01                   4
DME-OO                  C   2H   5O   3     G    300.00   3500.00 1800.00      1
 1.28946547e+01 1.03828282e-02-3.02554576e-06 3.64875471e-10-1.24113546e-14    2
-2.39005733e+04-3.76069562e+01 3.24067828e+00 3.18361092e-02-2.09032799e-05    3
 6.98625850e-09-9.32047886e-13-2.04251417e+04 1.46423783e+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   3500.00 1250.00      1
 1.07374983e+01 1.39769747e-02-5.32012597e-06 9.94916579e-10-7.50061107e-14    2
-1.73025108e+04-2.35990435e+01 1.12063956e-01 4.79783646e-02-4.61217939e-05    3
 2.27558061e-08-4.42718402e-12-1.46461523e+04 3.00335324e+01                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   3500.00 1370.00      1
 1.59411121e+01 1.44932690e-02-5.65697248e-06 1.09027852e-09-8.49010939e-14    2
-3.74943649e+04-4.65328702e+01 2.39014311e+00 5.40581418e-02-4.89761763e-05    3
 2.21701831e-08-3.93159900e-12-3.37813994e+04 2.31087123e+01                   4
DME-OQOOH               C   2H   4O   4     G    300.00   3500.00 1760.00      1
 1.54960865e+01 1.58758105e-03 2.24425902e-06-9.74237208e-10 1.03773066e-13    2
-4.69655432e+04-5.18401165e+01 3.62388957e+00 2.85698467e-02-2.07519902e-05    3
 7.73646324e-09-1.13354234e-12-4.27865299e+04 1.21478877e+01                   4
MTBE                    C   5H  12O   1     G    300.00   3500.00 1320.00      1
 9.85250856e+00 4.01896195e-02-1.66704212e-05 3.10158952e-09-2.11537798e-13    2
-4.09274217e+04-2.61941110e+01-1.85856423e+00 7.56777188e-02-5.69978069e-05    3
 2.34689560e-08-4.06899357e-12-3.78356985e+04 3.35564111e+01                   4
ETBE                    C   6H  14O   1     G    300.00   3500.00 1280.00      1
 1.16559136e+01 4.67933986e-02-1.93342013e-05 3.59185139e-09-2.45564974e-13    2
-4.60322114e+04-3.38084940e+01-3.48005605e+00 9.40933039e-02-7.47637779e-05    3
 3.24614225e-08-5.88415308e-12-4.21574031e+04 4.29502771e+01                   4
DIPE                    C   6H  14O   1     G    300.00   3500.00 1380.00      1
 1.11573928e+01 4.99175658e-02-2.25561386e-05 4.38444843e-09-3.06549364e-13    2
-4.59357929e+04-3.06117764e+01-2.50745274e+00 8.95258138e-02-6.56085821e-05    3
 2.51827303e-08-4.07435405e-12-4.21642955e+04 3.97144256e+01                   4
TAME                    C   6H  14O   1     G    300.00   3500.00 1320.00      1
 1.13309761e+01 4.74280943e-02-1.96957502e-05 3.66860749e-09-2.50688227e-13    2
-4.42745214e+04-3.17952395e+01-2.12836721e+00 8.82139832e-02-6.60433512e-05    3
 2.70764868e-08-4.68399870e-12-4.07212548e+04 3.68750527e+01                   4
RMTBE                   C   5H  11O   1     G    300.00   3500.00 1370.00      1
 1.09269229e+01 3.74766265e-02-1.73062474e-05 3.86241413e-09-3.39119740e-13    2
-1.88007827e+04-2.53563680e+01-1.81069451e-01 6.99087211e-02-5.28158399e-05    3
 2.11420212e-08-3.49233271e-12-1.57571928e+04 3.17301895e+01                   4
RDIPE                   C   6H  13O   1     G    300.00   3500.00 1800.00      1
 1.69549494e+01 3.45118423e-02-1.31342732e-05 2.36150212e-09-1.67133125e-13    2
-2.78147477e+04-5.54607976e+01 6.91787207e-01 7.06522027e-02-4.32512401e-05    3
 1.35159343e-08-1.71635982e-12-2.19600093e+04 3.25588287e+01                   4
MTBE-O                  C   5H  10O   2     G    300.00   3500.00 1520.00      1
 1.51388759e+01 2.99979380e-02-1.22799224e-05 2.46100800e-09-1.97690795e-13    2
-5.39879921e+04-5.57113238e+01-5.03717524e+00 8.30928094e-02-6.46761770e-05    3
 2.54418214e-08-3.97742985e-12-4.78544725e+04 5.00743811e+01                   4
MTBE-OO                 C   5H  11O   3     G    300.00   3500.00 1650.00      1
 1.64806404e+01 3.48147986e-02-1.47688716e-05 3.00165535e-09-2.41352124e-13    2
-3.59678540e+04-5.02874924e+01 2.84930352e+00 6.78604638e-02-4.48103854e-05    3
 1.51396407e-08-2.08044082e-12-3.14695128e+04 2.23020650e+01                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   3500.00 1320.00      1
 1.54436171e+01 3.66620452e-02-1.53964703e-05 3.18866664e-09-2.64826209e-13    2
-2.86187067e+04-4.25445321e+01 1.39866728e+00 7.92224991e-02-6.37606224e-05    3
 2.76150061e-08-4.89102686e-12-2.49108399e+04 2.91135557e+01                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   3500.00 1360.00      1
 1.70053287e+01 4.31260455e-02-1.99573148e-05 4.44658587e-09-3.89314848e-13    2
-4.64302952e+04-4.61328184e+01 4.65469152e+00 7.94514489e-02-6.00220979e-05    3
 2.40861854e-08-3.99953535e-12-4.30709219e+04 1.72494984e+01                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   3500.00 1750.00      1
 2.60727575e+01 2.16561734e-02-7.50837023e-06 1.18094191e-09-6.95946676e-14    2
-6.60762157e+04-1.03020582e+02 2.39248713e+00 7.57825058e-02-5.39023694e-05    3
 1.88548464e-08-2.59443816e-12-5.77881211e+04 2.44748876e+01                   4
CSOLID                  C   1               G    300.00   4000.00 1000.00      1
 .159828070E+01 .143065097E-02-.509435105E-06 .864401302E-10-.534349530E-14    2
-.745940284E+03-.930332005E+01-.303744539E+00 .436036227E-02 .198268825E-05    3
-.643472598E-08 .299601320E-11-.109458288E+03 .108301475E+01                   4
BIN1A                   C  20H  16          G   300.00   4000.00  1000.00      1
 .384004130e+02 .613760802e-01-.226838420e-04 .377828116e-08-.235041851e-12    2
-.165747108e+04-.190858878e+03-.946290891e+01 .179252381e+00-.989756752e-04    3
-.116559979e-07 .214782048e-10 .122142317e+05 .597553003e+02                   4
BIN1B                   C  20H  10          G   300.00   4000.00  1000.00      1
 .329670254e+02 .526917977e-01-.194742383e-04 .324368101e-08-.201785086e-12    2
 .107718330e+04-.161481167e+03-.895697031e+01 .146820540e+00-.577692501e-04    3
-.392441219e-07 .283752285e-10 .136083600e+05 .601566475e+02                   4
BIN1C                   C  20H   5          G   300.00   4000.00  1000.00      1
 .288518394e+02 .461144212e-01-.170433212e-04 .283878100e-08-.176596796e-12    2
-.612310898e+04-.152441597e+03-.829114243e+01 .126981825e+00-.389276128e-04    3
-.485387475e-07 .293596977e-10 .481805809e+04 .439495435e+02                   4
BIN2A                   C  40H  31          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .397395323e+03-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .283409758e+05 .136281912e+03                   4
BIN2B                   C  40H  16          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
-.435148944e+04-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .195176885e+05 .109755604e+03                   4
BIN2C                   C  40H   8          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
-.170085815e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .447424565e+04 .886402226e+02                   4
BIN3A                   C  80H  60          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .303189596e+04-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .578481001e+05 .254746237e+03                   4
BIN3B                   C  80H  24          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
-.213600710e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .239919342e+05 .198395827e+03                   4
BIN3C                   C  80H   8          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
-.466742552e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09-.609495158e+04 .156165064e+03                   4
BIN4A                   C 160H 116          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .105380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .118028497e+06 .473857298e+03                   4
BIN4B                   C 160H  32          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.680343262e+05-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .178969826e+05 .354560890e+03                   4
BIN4C                   C 160H  10          G   300.00   4000.00  1000.00      1
 .205435737e+03 .328351689e+00-.121354734e-03 .202131681e-07-.125743435e-11    2
-.102752674e+06-.113842566e+04-.653585808e+02 .890818250e+00-.172909327e-03    3
-.471736610e-06 .250565077e-09-.233838303e+05 .296493591e+03                   4
BIN5Aliq                C 320H 224          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .352119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .247380465e+06 .927804457e+03                   4
BIN5Bliq                C 320H  64          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.135714032e+06-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .361485852e+05 .709121781e+03                   4
BIN5Cliq                C 320H  18          G   300.00   4000.00  1000.00      1
 .409205747e+03 .654041015e+00-.241725492e-03 .402624424e-07-.250467310e-11    2
-.208758277e+06-.227246778e+04-.130537242e+03 .177352947e+01-.337554521e-03    3
-.947981323e-06 .501803389e-09-.506171764e+05 .587708337e+03                   4
BIN6Aliq                C 640H 432          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .909146192e+05-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .507419557e+06 .173874832e+04                   4
BIN6Bliq                C 640H 128          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.271428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .722971705e+05 .141824356e+04                   4
BIN6Cliq                C 640H  34          G   300.00   4000.00  1000.00      1
 .816745766e+03 .130541967e+01-.482467007e-03 .803609911e-07-.499915059e-11    2
-.420769482e+06-.454055202e+04-.260894565e+03 .353895191e+01-.666844909e-03    3
-.190047075e-05 .100428001e-08-.105083869e+06 .117013783e+04                   4
BIN7Aliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          813
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .219703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .101891965e+07 .319868647e+04                   4
BIN7Bliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          250
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.528501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .142639667e+06 .276398698e+04                   4
BIN7Cliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           65
 .159398623e+04 .254769728e+01-.941597491e-03 .156834989e-06-.975649647e-11    2
-.824746508e+06-.886326423e+04-.509649220e+03 .690588633e+01-.129480205e-02    3
-.371700233e-05 .196265639e-08-.208493980e+06 .228472375e+04                   4
BIN8Aliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1563
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .525439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .209454960e+07 .599019956e+04                   4
BIN8Bliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          500
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.106037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .282300003e+06 .554001391e+04                   4
BIN8Cliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          126
 .318473927e+04 .509022690e+01-.188128508e-02 .313351859e-06-.194932032e-10    2
-.165413482e+07-.177215999e+05-.101850654e+04 .137964163e+02-.257671322e-02    3
-.743906960e-05 .392526201e-08-.423020017e+06 .455286982e+04                   4
BIN9A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         3000
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .105415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .433609933e+07 .163588732e+05                   4
BIN9Aliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         3000
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .105415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .433609933e+07 .163588732e+05                   4
BIN9B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         1000
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.212075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .564600007e+06 .110800278e+05                   4
BIN9Bliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         1000
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.212075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .564600007e+06 .110800278e+05                   4
BIN9C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          251
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.330896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.847131304e+06 .910009023e+04                   4
BIN9Cliq                C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          251
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.330896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.847131304e+06 .910009023e+04                   4
BIN10A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5750
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .171313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .820225091e+07 .320518708e+05                   4
BIN10Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5750
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .171313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .820225091e+07 .320518708e+05                   4
BIN10AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5750
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .171313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .820225091e+07 .320518708e+05                   4
BIN10B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         2000
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.424150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .112920001e+07 .221600556e+05                   4
BIN10Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         2000
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.424150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .112920001e+07 .221600556e+05                   4
BIN10BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         2000
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.424150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .112920001e+07 .221600556e+05                   4
BIN10C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          501
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.662199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.169833321e+07 .182065710e+05                   4
BIN10Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          501
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.662199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.169833321e+07 .182065710e+05                   4
BIN10CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          501
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.662199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.169833321e+07 .182065710e+05                   4
BIN11A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        11000
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .262917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .154586477e+08 .627960702e+05                   4
BIN11Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        11000
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .262917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .154586477e+08 .627960702e+05                   4
BIN11AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        11000
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .262917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .154586477e+08 .627960702e+05                   4
BIN11B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         4000
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.848301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .225840003e+07 .443201113e+05                   4
BIN11Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         4000
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.848301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .225840003e+07 .443201113e+05                   4
BIN11BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         4000
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.848301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .225840003e+07 .443201113e+05                   4
BIN11C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1001
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.132446866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.339775769e+07 .364074926e+05                   4
BIN11Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1001
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.132446866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.339775769e+07 .364074926e+05                   4
BIN11CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1001
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.132446866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.339775769e+07 .364074926e+05                   4
BIN12A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        21000
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .367089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290315457e+08 .122952718e+06                   4
BIN12Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        21000
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .367089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290315457e+08 .122952718e+06                   4
BIN12AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        21000
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .367089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290315457e+08 .122952718e+06                   4
BIN12B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         8000
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169660271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .451680005e+07 .886402226e+05                   4
BIN12Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         8000
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169660271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .451680005e+07 .886402226e+05                   4
BIN12BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         8000
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169660271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .451680005e+07 .886402226e+05                   4
BIN12C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2001
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264900676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.679660664e+07 .728093358e+05                   4
BIN12Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2001
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264900676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.679660664e+07 .728093358e+05                   4
BIN12CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2001
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264900676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.679660664e+07 .728093358e+05                   4
BIN13A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        40000
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .416688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .542915920e+08 .240626590e+06                   4
BIN13Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        40000
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .416688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .542915920e+08 .240626590e+06                   4
BIN13AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        40000
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .416688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .542915920e+08 .240626590e+06                   4
BIN13B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        16000
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.339320543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .903360011e+07 .177280445e+06                   4
BIN13Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        16000
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.339320543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .903360011e+07 .177280445e+06                   4
BIN13BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        16000
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.339320543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .903360011e+07 .177280445e+06                   4
BIN13C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4001
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529808296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135943046e+08 .145613022e+06                   4
BIN13Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4001
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529808296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135943046e+08 .145613022e+06                   4
BIN13CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4001
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529808296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135943046e+08 .145613022e+06                   4
BIN14A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        76000
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .198394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101040185e+09 .470695489e+06                   4
BIN14Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        76000
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .198394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101040185e+09 .470695489e+06                   4
BIN14AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        76000
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .198394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101040185e+09 .470695489e+06                   4
BIN14B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        32000
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678641086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .180672002e+08 .354560890e+06                   4
BIN14Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        32000
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678641086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .180672002e+08 .354560890e+06                   4
BIN14BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        32000
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678641086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .180672002e+08 .354560890e+06                   4
BIN14C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8001
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105962354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271897004e+08 .291220395e+06                   4
BIN14Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8001
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105962354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271897004e+08 .291220395e+06                   4
BIN14CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8001
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105962354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271897004e+08 .291220395e+06                   4
BIN15A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       144000
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.873175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .186994373e+09 .920275597e+06                   4
BIN15Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       144000
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.873175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .186994373e+09 .920275597e+06                   4
BIN15AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       144000
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.873175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .186994373e+09 .920275597e+06                   4
BIN15B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        64000
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135728217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361344004e+08 .709121781e+06                   4
BIN15Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        64000
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135728217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361344004e+08 .709121781e+06                   4
BIN15BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        64000
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135728217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361344004e+08 .709121781e+06                   4
BIN15C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16001
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211925402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543804920e+08 .582435141e+06                   4
BIN15Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16001
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211925402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543804920e+08 .582435141e+06                   4
BIN15CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16001
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211925402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543804920e+08 .582435141e+06                   4
BIN16A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32001
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423851498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108762075e+09 .116486463e+07                   4
BIN16Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32001
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423851498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108762075e+09 .116486463e+07                   4
BIN16CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32001
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423851498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108762075e+09 .116486463e+07                   4
BIN16CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32001
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423851498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108762075e+09 .116486463e+07                   4
BIN17A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       512000
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136524181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627289515e+09 .351217933e+07                   4
BIN17Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       512000
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136524181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627289515e+09 .351217933e+07                   4
BIN17AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       512000
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136524181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627289515e+09 .351217933e+07                   4
BIN17AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       512000
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136524181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627289515e+09 .351217933e+07                   4
BIN17B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       256000
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542912868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144537602e+09 .283648712e+07                   4
BIN17Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       256000
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542912868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144537602e+09 .283648712e+07                   4
BIN17BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       256000
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542912868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144537602e+09 .283648712e+07                   4
BIN17BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       256000
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542912868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144537602e+09 .283648712e+07                   4
BIN17C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64001
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847703690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217525242e+09 .232972361e+07                   4
BIN17Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64001
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847703690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217525242e+09 .232972361e+07                   4
BIN17CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64001
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847703690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217525242e+09 .232972361e+07                   4
BIN17CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64001
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847703690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217525242e+09 .232972361e+07                   4
BIN18A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       960000
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374645533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113389105e+10 .685543562e+07                   4
BIN18Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       960000
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374645533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113389105e+10 .685543562e+07                   4
BIN18AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       960000
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374645533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113389105e+10 .685543562e+07                   4
BIN18AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       960000
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374645533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113389105e+10 .685543562e+07                   4
BIN18B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       512000
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108582574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289075203e+09 .567297425e+07                   4
BIN18Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       512000
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108582574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289075203e+09 .567297425e+07                   4
BIN18BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       512000
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108582574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289075203e+09 .567297425e+07                   4
BIN18BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       512000
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108582574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289075203e+09 .567297425e+07                   4
BIN18C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128001
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169540807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.435051575e+09 .465944158e+07                   4
BIN18Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128001
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169540807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.435051575e+09 .465944158e+07                   4
BIN18CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128001
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169540807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.435051575e+09 .465944158e+07                   4
BIN18CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128001
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169540807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.435051575e+09 .465944158e+07                   4
BIN19A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1792000
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952485410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202640615e+10 .133730251e+08                   4
BIN19Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1792000
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952485410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202640615e+10 .133730251e+08                   4
BIN19AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1792000
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952485410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202640615e+10 .133730251e+08                   4
BIN19AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1792000
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952485410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202640615e+10 .133730251e+08                   4
BIN19B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1024000
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217165147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578150407e+09 .113459485e+08                   4
BIN19Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1024000
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217165147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578150407e+09 .113459485e+08                   4
BIN19BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1024000
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217165147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578150407e+09 .113459485e+08                   4
BIN19BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1024000
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217165147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578150407e+09 .113459485e+08                   4
BIN19C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256001
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339081684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870104242e+09 .931887751e+07                   4
BIN19Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256001
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339081684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870104242e+09 .931887751e+07                   4
BIN19CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256001
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339081684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870104242e+09 .931887751e+07                   4
BIN19CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256001
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339081684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870104242e+09 .931887751e+07                   4
BIN20A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3328000
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231135951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357006038e+10 .260703580e+08                   4
BIN20Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3328000
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231135951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357006038e+10 .260703580e+08                   4
BIN20AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3328000
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231135951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357006038e+10 .260703580e+08                   4
BIN20AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3328000
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231135951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357006038e+10 .260703580e+08                   4
BIN20B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2048000
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434330295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115630081e+10 .226918970e+08                   4
BIN20Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2048000
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434330295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115630081e+10 .226918970e+08                   4
BIN20BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2048000
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434330295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115630081e+10 .226918970e+08                   4
BIN20BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2048000
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434330295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115630081e+10 .226918970e+08                   4
BIN20C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512001
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678163438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174020957e+10 .186377494e+08                   4
BIN20Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512001
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678163438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174020957e+10 .186377494e+08                   4
BIN20CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512001
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678163438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174020957e+10 .186377494e+08                   4
BIN20CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512001
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678163438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174020957e+10 .186377494e+08                   4
BIN21A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6144000
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543549639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617461693e+10 .507893317e+08                   4
BIN21Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6144000
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543549639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617461693e+10 .507893317e+08                   4
BIN21AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6144000
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543549639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617461693e+10 .507893317e+08                   4
BIN21AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6144000
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543549639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617461693e+10 .507893317e+08                   4
BIN21B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4096000
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868660590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231260163e+10 .453837940e+08                   4
BIN21Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4096000
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868660590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231260163e+10 .453837940e+08                   4
BIN21BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4096000
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868660590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231260163e+10 .453837940e+08                   4
BIN21BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4096000
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868660590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231260163e+10 .453837940e+08                   4
BIN21C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024001
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632695e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348042024e+10 .372754931e+08                   4
BIN21Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024001
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632695e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348042024e+10 .372754931e+08                   4
BIN21CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024001
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632695e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348042024e+10 .372754931e+08                   4
BIN21CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024001
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632695e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348042024e+10 .372754931e+08                   4
BIN22A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12288000
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709928e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492339e+11 .101578663e+09                   4
BIN22Aliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12288000
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709928e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492339e+11 .101578663e+09                   4
BIN22AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12288000
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709928e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492339e+11 .101578663e+09                   4
BIN22AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12288000
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709928e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492339e+11 .101578663e+09                   4
BIN22B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8192000
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173732118e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462520326e+10 .907675879e+08                   4
BIN22Bliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8192000
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173732118e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462520326e+10 .907675879e+08                   4
BIN22BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8192000
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173732118e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462520326e+10 .907675879e+08                   4
BIN22BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8192000
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173732118e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462520326e+10 .907675879e+08                   4
BIN22C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048001
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271265403e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696084266e+10 .745509749e+08                   4
BIN22Cliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048001
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271265403e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696084266e+10 .745509749e+08                   4
BIN22CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048001
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271265403e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696084266e+10 .745509749e+08                   4
BIN22CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048001
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271265403e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696084266e+10 .745509749e+08                   4
BIN23AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24576000
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419856e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246984677e+11 .203157327e+09                   4
BIN23AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24576000
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419856e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246984677e+11 .203157327e+09                   4
BIN23AaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24576000
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419856e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246984677e+11 .203157327e+09                   4
BIN23BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16384000
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347464236e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925040651e+10 .181535176e+09                   4
BIN23BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16384000
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347464236e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925040651e+10 .181535176e+09                   4
BIN23BaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16384000
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347464236e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925040651e+10 .181535176e+09                   4
BIN23CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096001
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530799e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216842e+11 .149101955e+09                   4
BIN23CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096001
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530799e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216842e+11 .149101955e+09                   4
BIN23CaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096001
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530799e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216842e+11 .149101955e+09                   4
BIN24AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49152000
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839711e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969355e+11 .406314653e+09                   4
BIN24AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49152000
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839711e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969355e+11 .406314653e+09                   4
BIN24AaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49152000
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839711e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969355e+11 .406314653e+09                   4
BIN24BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32768000
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694928472e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008130e+11 .363070352e+09                   4
BIN24BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32768000
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694928472e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008130e+11 .363070352e+09                   4
BIN24BaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32768000
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694928472e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008130e+11 .363070352e+09                   4
BIN24CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192001
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506160e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433696e+11 .298203905e+09                   4
BIN24CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192001
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506160e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433696e+11 .298203905e+09                   4
BIN24CaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192001
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506160e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433696e+11 .298203905e+09                   4
BIN25AaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98304000
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869679423e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987938710e+11 .812629307e+09                   4
BIN25AaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98304000
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869679423e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987938710e+11 .812629307e+09                   4
BIN25AaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98304000
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869679423e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987938710e+11 .812629307e+09                   4
BIN25BaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65536000
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985694e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016260e+11 .726140704e+09                   4
BIN25BaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65536000
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985694e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016260e+11 .726140704e+09                   4
BIN25BaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65536000
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985694e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016260e+11 .726140704e+09                   4
BIN25CaggI              C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384001
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012322e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556867402e+11 .596407805e+09                   4
BIN25CaggII             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384001
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012322e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556867402e+11 .596407805e+09                   4
BIN25CaggIII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384001
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012322e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556867402e+11 .596407805e+09                   4
BIN1AJ                  C  20H  15          G   300.00   4000.00  1000.00      1
 .384004130e+02 .613760802e-01-.226838420e-04 .377828116e-08-.235041851e-12    2
 .583425289e+05-.190858878e+03-.946290891e+01 .179252381e+00-.989756752e-04    3
-.116559979e-07 .214782048e-10 .722142317e+05 .597553003e+02                   4
BIN1BJ                  C  20H   9          G   300.00   4000.00  1000.00      1
 .329670254e+02 .526917977e-01-.194742383e-04 .324368101e-08-.201785086e-12    2
 .610771833e+05-.161481167e+03-.895697031e+01 .146820540e+00-.577692501e-04    3
-.392441219e-07 .283752285e-10 .736083600e+05 .601566475e+02                   4
BIN1CJ                  C  20H   4          G   300.00   4000.00  1000.00      1
 .288518394e+02 .461144212e-01-.170433212e-04 .283878100e-08-.176596796e-12    2
 .538768910e+05-.152441597e+03-.829114243e+01 .126981825e+00-.389276128e-04    3
-.485387475e-07 .293596977e-10 .648180581e+05 .439495435e+02                   4
BIN2AJ                  C  40H  30          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .603973953e+05-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .883409758e+05 .136281912e+03                   4
BIN2BJ                  C  40H  15          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
 .556485106e+05-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .795176885e+05 .109755604e+03                   4
BIN2CJ                  C  40H   7          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
 .429914185e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .644742457e+05 .886402226e+02                   4
BIN3AJ                  C  80H  59          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .630318960e+05-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .117848100e+06 .254746237e+03                   4
BIN3BJ                  C  80H  23          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
 .386399290e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .839919342e+05 .198395827e+03                   4
BIN3CJ                  C  80H   7          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
 .133257448e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09 .539050484e+05 .156165064e+03                   4
BIN4AJ                  C 160H 115          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .705380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .178028497e+06 .473857298e+03                   4
BIN4BJ                  C 160H  31          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.803432616e+04-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .778969826e+05 .354560890e+03                   4
BIN4CJ                  C 160H   9          G   300.00   4000.00  1000.00      1
 .205435737e+03 .328351689e+00-.121354734e-03 .202131681e-07-.125743435e-11    2
-.427526744e+05-.113842566e+04-.653585808e+02 .890818250e+00-.172909327e-03    3
-.471736610e-06 .250565077e-09 .366161697e+05 .296493591e+03                   4
BIN5AJliq               C 320H 223          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .952119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .307380465e+06 .927804457e+03                   4
BIN5BJliq               C 320H  63          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.757140323e+05-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .961485852e+05 .709121781e+03                   4
BIN5CJliq               C 320H  17          G   300.00   4000.00  1000.00      1
 .409205747e+03 .654041015e+00-.241725492e-03 .402624424e-07-.250467310e-11    2
-.148758277e+06-.227246778e+04-.130537242e+03 .177352947e+01-.337554521e-03    3
-.947981323e-06 .501803389e-09 .938282361e+04 .587708337e+03                   4
BIN6AJliq               C 640H 431          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .150914619e+06-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .567419557e+06 .173874832e+04                   4
BIN6BJliq               C 640H 127          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.211428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .132297170e+06 .141824356e+04                   4
BIN6CJliq               C 640H  33          G   300.00   4000.00  1000.00      1
 .816745766e+03 .130541967e+01-.482467007e-03 .803609911e-07-.499915059e-11    2
-.360769482e+06-.454055202e+04-.260894565e+03 .353895191e+01-.666844909e-03    3
-.190047075e-05 .100428001e-08-.450838685e+05 .117013783e+04                   4
BIN7AJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          812
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .279703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .107891965e+07 .319868647e+04                   4
BIN7BJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          249
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.468501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .202639667e+06 .276398698e+04                   4
BIN7CJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           64
 .159398623e+04 .254769728e+01-.941597491e-03 .156834989e-06-.975649647e-11    2
-.764746508e+06-.886326423e+04-.509649220e+03 .690588633e+01-.129480205e-02    3
-.371700233e-05 .196265639e-08-.148493980e+06 .228472375e+04                   4
BIN8AJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1562
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .585439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .215454960e+07 .599019956e+04                   4
BIN8BJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          499
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.100037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .342300003e+06 .554001391e+04                   4
BIN8CJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          125
 .318473927e+04 .509022690e+01-.188128508e-02 .313351859e-06-.194932032e-10    2
-.159413482e+07-.177215999e+05-.101850654e+04 .137964163e+02-.257671322e-02    3
-.743906960e-05 .392526201e-08-.363020017e+06 .455286982e+04                   4
BIN9AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         2999
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .111415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .439609933e+07 .163588732e+05                   4
BIN9AJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         2999
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .111415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .439609933e+07 .163588732e+05                   4
BIN9BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          999
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.206075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .624600007e+06 .110800278e+05                   4
BIN9BJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          999
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.206075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .624600007e+06 .110800278e+05                   4
BIN9CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          250
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.324896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.787131304e+06 .910009023e+04                   4
BIN9CJliq               C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          250
 .636869480e+04 .101792011e+02-.376210719e-02 .626626605e-06-.389816093e-10    2
-.324896407e+07-.354429274e+05-.203670710e+04 .275892080e+02-.515111307e-02    3
-.148784176e-04 .785016202e-08-.787131304e+06 .910009023e+04                   4
BIN10AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5749
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .177313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .826225091e+07 .320518708e+05                   4
BIN10AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5749
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .177313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .826225091e+07 .320518708e+05                   4
BIN10AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5749
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .177313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .826225091e+07 .320518708e+05                   4
BIN10BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         1999
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.418150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .118920001e+07 .221600556e+05                   4
BIN10BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         1999
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.418150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .118920001e+07 .221600556e+05                   4
BIN10BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         1999
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.418150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .118920001e+07 .221600556e+05                   4
BIN10CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          500
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.656199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.163833321e+07 .182065710e+05                   4
BIN10CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          500
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.656199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.163833321e+07 .182065710e+05                   4
BIN10CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          500
 .127364093e+05 .203568355e+02-.752363532e-02 .125315676e-05-.779572186e-10    2
-.656199607e+07-.708779052e+05-.407397232e+04 .551730759e+02-.102926380e-01    3
-.297650162e-04 .157027565e-07-.163833321e+07 .182065710e+05                   4
BIN11AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        10999
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .268917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .155186477e+08 .627960702e+05                   4
BIN11AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        10999
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .268917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .155186477e+08 .627960702e+05                   4
BIN11AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        10999
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .268917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .155186477e+08 .627960702e+05                   4
BIN11BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         3999
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.842301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .231840003e+07 .443201113e+05                   4
BIN11BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         3999
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.842301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .231840003e+07 .443201113e+05                   4
BIN11BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         3999
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.842301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .231840003e+07 .443201113e+05                   4
BIN11CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1000
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.131846866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.333775769e+07 .364074926e+05                   4
BIN11CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1000
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.131846866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.333775769e+07 .364074926e+05                   4
BIN11CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1000
 .254720349e+05 .407124184e+02-.150468077e-01 .250623641e-05-.155909640e-09    2
-.131846866e+08-.141755538e+06-.814763865e+04 .110342527e+03-.205829626e-01    3
-.595303108e-04 .314051510e-07-.333775769e+07 .364074926e+05                   4
BIN12AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        20999
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .373089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290915457e+08 .122952718e+06                   4
BIN12AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        20999
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .373089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290915457e+08 .122952718e+06                   4
BIN12AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        20999
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .373089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290915457e+08 .122952718e+06                   4
BIN12BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         7999
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169060271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .457680005e+07 .886402226e+05                   4
BIN12BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         7999
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169060271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .457680005e+07 .886402226e+05                   4
BIN12BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         7999
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169060271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .457680005e+07 .886402226e+05                   4
BIN12CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2000
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264300676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.673660664e+07 .728093358e+05                   4
BIN12CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2000
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264300676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.673660664e+07 .728093358e+05                   4
BIN12CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2000
 .509432862e+05 .814235841e+02-.300931524e-01 .501239570e-05-.311814483e-09    2
-.264300676e+08-.283510803e+06-.162949713e+05 .220681430e+03-.411636118e-01    3
-.119060900e-03 .628099400e-07-.673660664e+07 .728093358e+05                   4
BIN13AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        39999
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .422688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .543515920e+08 .240626590e+06                   4
BIN13AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        39999
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .422688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .543515920e+08 .240626590e+06                   4
BIN13AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        39999
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .422688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .543515920e+08 .240626590e+06                   4
BIN13BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        15999
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.338720543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .909360011e+07 .177280445e+06                   4
BIN13BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        15999
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.338720543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .909360011e+07 .177280445e+06                   4
BIN13BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        15999
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.338720543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .909360011e+07 .177280445e+06                   4
BIN13CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4000
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529208296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135343046e+08 .145613022e+06                   4
BIN13CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4000
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529208296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135343046e+08 .145613022e+06                   4
BIN13CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4000
 .101885789e+06 .162845916e+03-.601858418e-01 .100247143e-04-.623624169e-09    2
-.529208296e+08-.567021334e+06-.325896366e+05 .441359234e+03-.823249102e-01    3
-.238122078e-03 .125619518e-06-.135343046e+08 .145613022e+06                   4
BIN14AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        75999
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .204394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101100185e+09 .470695489e+06                   4
BIN14AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        75999
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .204394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101100185e+09 .470695489e+06                   4
BIN14AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        75999
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .204394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101100185e+09 .470695489e+06                   4
BIN14BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        31999
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678041086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .181272002e+08 .354560890e+06                   4
BIN14BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        31999
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678041086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .181272002e+08 .354560890e+06                   4
BIN14BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        31999
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678041086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .181272002e+08 .354560890e+06                   4
BIN14CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8000
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105902354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271297004e+08 .291220395e+06                   4
BIN14CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8000
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105902354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271297004e+08 .291220395e+06                   4
BIN14CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8000
 .203770793e+06 .325690579e+03-.120371221e+00 .200493515e-04-.124724354e-08    2
-.105902354e+09-.113404239e+07-.651789673e+05 .882714844e+03-.164647507e+00    3
-.476244435e-03 .251238674e-06-.271297004e+08 .291220395e+06                   4
BIN15AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       143999
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.867175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .187054373e+09 .920275597e+06                   4
BIN15AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       143999
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.867175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .187054373e+09 .920275597e+06                   4
BIN15AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       143999
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.867175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .187054373e+09 .920275597e+06                   4
BIN15BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        63999
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135668217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361944004e+08 .709121781e+06                   4
BIN15BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        63999
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135668217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361944004e+08 .709121781e+06                   4
BIN15BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        63999
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135668217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361944004e+08 .709121781e+06                   4
BIN15CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16000
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211865402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543204920e+08 .582435141e+06                   4
BIN15CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16000
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211865402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543204920e+08 .582435141e+06                   4
BIN15CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16000
 .407540803e+06 .651379905e+03-.240741978e+00 .400986258e-04-.249448229e-08    2
-.211865402e+09-.226808452e+07-.130357629e+06 .176542606e+04-.329292701e+00    3
-.952489148e-03 .502476986e-06-.543204920e+08 .582435141e+06                   4
BIN16AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423791498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108702075e+09 .116486463e+07                   4
BIN16CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423791498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108702075e+09 .116486463e+07                   4
BIN16CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423791498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108702075e+09 .116486463e+07                   4
BIN16CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080823e+06 .130275856e+04-.481483494e+00 .801971745e-04-.498895977e-08    2
-.423791498e+09-.453616876e+07-.260714951e+06 .353084850e+04-.658583088e+00    3
-.190497858e-02 .100495361e-05-.108702075e+09 .116486463e+07                   4
BIN17AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       511999
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136464181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627349515e+09 .351217933e+07                   4
BIN17AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       511999
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136464181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627349515e+09 .351217933e+07                   4
BIN17AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       511999
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136464181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627349515e+09 .351217933e+07                   4
BIN17AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       511999
 .200328306e+07 .320188384e+04-.118337677e+01 .197106387e-03-.122617265e-07    2
-.136464181e+09-.100542485e+08-.561731253e+06 .887766459e+04-.316832746e+01    3
-.280014245e-02 .185910170e-05 .627349515e+09 .351217933e+07                   4
BIN17BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       255999
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542852868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144597602e+09 .283648712e+07                   4
BIN17BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       255999
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542852868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144597602e+09 .283648712e+07                   4
BIN17BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       255999
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542852868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144597602e+09 .283648712e+07                   4
BIN17BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H       255999
 .179006993e+07 .286110142e+04-.105742779e+01 .176127992e-03-.109566885e-07    2
-.542852868e+09-.949315621e+07-.538701560e+06 .783996468e+04-.211051837e+01    3
-.337717974e-02 .194527587e-05 .144597602e+09 .283648712e+07                   4
BIN17CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64000
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847643690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217465242e+09 .232972361e+07                   4
BIN17CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64000
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847643690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217465242e+09 .232972361e+07                   4
BIN17CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64000
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847643690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217465242e+09 .232972361e+07                   4
BIN17CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      1280000 H        64000
 .163016086e+07 .260551586e+04-.962966525e+00 .160394272e-03-.997791475e-08    2
-.847643690e+09-.907233725e+07-.521429596e+06 .706169338e+04-.131716386e+01    3
-.380995743e-02 .200990686e-05-.217465242e+09 .232972361e+07                   4
BIN18AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       959999
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374585533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113395105e+10 .685543562e+07                   4
BIN18AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       959999
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374585533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113395105e+10 .685543562e+07                   4
BIN18AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       959999
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374585533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113395105e+10 .685543562e+07                   4
BIN18AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       959999
 .395326284e+07 .631857208e+04-.233526629e+01 .388968175e-03-.241971935e-07    2
-.374585533e+09-.199682240e+08-.111770508e+07 .174959042e+05-.607220265e+01    3
-.574454422e-02 .373974695e-05 .113395105e+10 .685543562e+07                   4
BIN18BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       511999
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108576574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289135203e+09 .567297425e+07                   4
BIN18BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       511999
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108576574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289135203e+09 .567297425e+07                   4
BIN18BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       511999
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108576574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289135203e+09 .567297425e+07                   4
BIN18BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       511999
 .358013985e+07 .572220284e+04-.211485558e+01 .352255983e-03-.219133769e-07    2
-.108576574e+10-.189863124e+08-.107740312e+07 .156799294e+05-.422103674e+01    3
-.675435948e-02 .389055174e-05 .289135203e+09 .567297425e+07                   4
BIN18CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128000
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169534807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.434991575e+09 .465944158e+07                   4
BIN18CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128000
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169534807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.434991575e+09 .465944158e+07                   4
BIN18CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128000
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169534807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.434991575e+09 .465944158e+07                   4
BIN18CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      2560000 H       128000
 .326032094e+07 .521103047e+04-.192593259e+01 .320788467e-03-.199558247e-07    2
-.169534807e+10-.181446742e+08-.104285889e+07 .141233831e+05-.263432541e+01    3
-.761991514e-02 .401981336e-05-.434991575e+09 .465944158e+07                   4
BIN19AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1791999
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952425410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202646615e+10 .133730251e+08                   4
BIN19AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1791999
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952425410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202646615e+10 .133730251e+08                   4
BIN19AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1791999
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952425410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202646615e+10 .133730251e+08                   4
BIN19AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1791999
 .779991911e+07 .124667529e+05-.460755809e+01 .767447153e-03-.477418679e-07    2
-.952425410e+09-.396559018e+08-.222389532e+07 .344729584e+05-.116155008e+02    3
-.117776071e-01 .752258099e-05 .202646615e+10 .133730251e+08                   4
BIN19BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1023999
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217159147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578210407e+09 .113459485e+08                   4
BIN19BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1023999
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217159147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578210407e+09 .113459485e+08                   4
BIN19BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1023999
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217159147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578210407e+09 .113459485e+08                   4
BIN19BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H      1023999
 .716027971e+07 .114444057e+05-.422971117e+01 .704511966e-03-.438267539e-07    2
-.217159147e+10-.379726248e+08-.215480624e+07 .313598587e+05-.844207348e+01    3
-.135087190e-01 .778110349e-05 .578210407e+09 .113459485e+08                   4
BIN19CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256000
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339075684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870044242e+09 .931887751e+07                   4
BIN19CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256000
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339075684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870044242e+09 .931887751e+07                   4
BIN19CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256000
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339075684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870044242e+09 .931887751e+07                   4
BIN19CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C      5120000 H       256000
 .652064109e+07 .104220597e+05-.385186471e+01 .641576856e-03-.399116446e-07    2
-.339075684e+10-.362893482e+08-.208571747e+07 .282467626e+05-.526864851e+01    3
-.152398306e-01 .803962635e-05-.870044242e+09 .931887751e+07                   4
BIN20AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3327999
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231129951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357012038e+10 .260703580e+08                   4
BIN20AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3327999
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231129951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357012038e+10 .260703580e+08                   4
BIN20AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3327999
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231129951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357012038e+10 .260703580e+08                   4
BIN20AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      3327999
 .153866251e+08 .245927235e+05-.908916721e+01 .151391591e-02-.941786978e-07    2
-.231129951e+10-.787507113e+08-.442476095e+07 .679082170e+05-.221731924e+02    3
-.241322514e-01 .151313361e-04 .357012038e+10 .260703580e+08                   4
BIN20BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2047999
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434324295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115636081e+10 .226918970e+08                   4
BIN20BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2047999
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434324295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115636081e+10 .226918970e+08                   4
BIN20BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2047999
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434324295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115636081e+10 .226918970e+08                   4
BIN20BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H      2047999
 .143205594e+08 .228888114e+05-.845942234e+01 .140902393e-02-.876535077e-07    2
-.434324295e+10-.759452497e+08-.430961248e+07 .627197175e+05-.168841470e+02    3
-.270174379e-01 .155622070e-04 .115636081e+10 .226918970e+08                   4
BIN20CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512000
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678157438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174014957e+10 .186377494e+08                   4
BIN20CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512000
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678157438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174014957e+10 .186377494e+08                   4
BIN20CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512000
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678157438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174014957e+10 .186377494e+08                   4
BIN20CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     10240000 H       512000
 .130412814e+08 .208441181e+05-.770372896e+01 .128315364e-02-.798232844e-07    2
-.678157438e+10-.725786961e+08-.417143463e+07 .564935217e+05-.105372947e+02    3
-.304796614e-01 .160792523e-04-.174014957e+10 .186377494e+08                   4
BIN21AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6143999
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543543639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617467693e+10 .507893317e+08                   4
BIN21AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6143999
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543543639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617467693e+10 .507893317e+08                   4
BIN21AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6143999
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543543639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617467693e+10 .507893317e+08                   4
BIN21AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      6143999
 .303468239e+08 .485038821e+05-.179264365e+02 .298587503e-02-.185747320e-06    2
-.543543639e+10-.156379238e+09-.880346251e+07 .133741034e+06-.422307666e+02    3
-.494185775e-01 .304350206e-04 .617467693e+10 .507893317e+08                   4
BIN21BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4095999
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868654590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231266163e+10 .453837940e+08                   4
BIN21BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4095999
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868654590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231266163e+10 .453837940e+08                   4
BIN21BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4095999
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868654590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231266163e+10 .453837940e+08                   4
BIN21BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      4095999
 .286411188e+08 .457776228e+05-.169188447e+02 .281804786e-02-.175307015e-06    2
-.868654590e+10-.151890499e+09-.861922496e+07 .125439435e+06-.337682939e+02    3
-.540348758e-01 .311244140e-04 .231266163e+10 .453837940e+08                   4
BIN21CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024000
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632095e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348036024e+10 .372754931e+08                   4
BIN21CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024000
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632095e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348036024e+10 .372754931e+08                   4
BIN21CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024000
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632095e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348036024e+10 .372754931e+08                   4
BIN21CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     20480000 H      1024000
 .260825620e+08 .416882350e+05-.154074575e+02 .256630719e-02-.159646564e-06    2
-.135632095e+11-.145157392e+09-.834286895e+07 .112987040e+06-.210745871e+02    3
-.609593230e-01 .321585043e-04-.348036024e+10 .372754931e+08                   4
BIN22AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12287999
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709328e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492939e+11 .101578663e+09                   4
BIN22AJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12287999
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709328e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492939e+11 .101578663e+09                   4
BIN22AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12287999
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709328e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492939e+11 .101578663e+09                   4
BIN22AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H     12287999
 .606936478e+08 .970077642e+05-.358528729e+02 .597175006e-02-.371494639e-06    2
-.108709328e+11-.312758476e+09-.176069250e+08 .267482068e+06-.844615333e+02    3
-.988371550e-01 .608700412e-04 .123492939e+11 .101578663e+09                   4
BIN22BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8191999
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173731518e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462526326e+10 .907675879e+08                   4
BIN22BJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8191999
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173731518e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462526326e+10 .907675879e+08                   4
BIN22BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8191999
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173731518e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462526326e+10 .907675879e+08                   4
BIN22BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      8191999
 .572822377e+08 .915552455e+05-.338376893e+02 .563609573e-02-.350614031e-06    2
-.173731518e+11-.303780999e+09-.172384499e+08 .250878870e+06-.675365878e+02    3
-.108069752e+00 .622488279e-04 .462526326e+10 .907675879e+08                   4
BIN22CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048000
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271264803e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696078266e+10 .745509749e+08                   4
BIN22CJliq              C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048000
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271264803e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696078266e+10 .745509749e+08                   4
BIN22CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048000
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271264803e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696078266e+10 .745509749e+08                   4
BIN22CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     40960000 H      2048000
 .521651225e+08 .833764675e+05-.308149140e+02 .513261423e-02-.319293119e-06    2
-.271264803e+11-.290314783e+09-.166857373e+08 .225974072e+06-.421491696e+02    3
-.121918647e+00 .643170079e-04-.696078266e+10 .745509749e+08                   4
BIN23AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24575999
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419256e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246985277e+11 .203157327e+09                   4
BIN23AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24575999
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419256e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246985277e+11 .203157327e+09                   4
BIN23AJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     24575999
 .121387296e+09 .194015528e+06-.717057459e+02 .119435001e-01-.742989279e-06    2
-.217419256e+11-.625516952e+09-.352138500e+08 .534964137e+06-.168923067e+03    3
-.197674310e+00 .121740082e-03 .246985277e+11 .203157327e+09                   4
BIN23BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16383999
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347463636e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925046651e+10 .181535176e+09                   4
BIN23BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16383999
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347463636e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925046651e+10 .181535176e+09                   4
BIN23BJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H     16383999
 .114564475e+09 .183110491e+06-.676753787e+02 .112721915e-01-.701228062e-06    2
-.347463636e+11-.607561998e+09-.344768998e+08 .501757740e+06-.135073176e+03    3
-.216139503e+00 .124497656e-03 .925046651e+10 .181535176e+09                   4
BIN23CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096000
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530199e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216242e+11 .149101955e+09                   4
BIN23CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096000
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530199e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216242e+11 .149101955e+09                   4
BIN23CJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C     81920000 H      4096000
 .104330246e+09 .166752936e+06-.616298284e+02 .102652285e-01-.638586242e-06    2
-.542530199e+11-.580629567e+09-.333714749e+08 .451948148e+06-.842983415e+02    3
-.243837293e+00 .128634016e-03-.139216242e+11 .149101955e+09                   4
BIN24AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49151999
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839111e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969955e+11 .406314653e+09                   4
BIN24AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49151999
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839111e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969955e+11 .406314653e+09                   4
BIN24AJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     49151999
 .242774591e+09 .388031057e+06-.143411492e+03 .238870002e-01-.148597856e-05    2
-.434839111e+11-.125103390e+10-.704277001e+08 .106992827e+07-.337846133e+03    3
-.395348620e+00 .243480165e-03 .493969955e+11 .406314653e+09                   4
BIN24BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32767999
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694927872e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008730e+11 .363070352e+09                   4
BIN24BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32767999
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694927872e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008730e+11 .363070352e+09                   4
BIN24BJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H     32767999
 .229128951e+09 .366220982e+06-.135350757e+03 .225443829e-01-.140245612e-05    2
-.694927872e+11-.121512400e+10-.689537997e+08 .100351548e+07-.270146351e+03    3
-.432279007e+00 .248995312e-03 .185008730e+11 .363070352e+09                   4
BIN24CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192000
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506100e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433096e+11 .298203905e+09                   4
BIN24CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192000
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506100e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433096e+11 .298203905e+09                   4
BIN24CJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    163840000 H      8192000
 .208660491e+09 .333505871e+06-.123259656e+03 .205304570e-01-.127717248e-05    2
-.108506100e+12-.116125913e+10-.667429495e+08 .903896292e+06-.168596681e+03    3
-.487674586e+00 .257268032e-03-.278433096e+11 .298203905e+09                   4
BIN25AJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98303999
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869678823e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987939310e+11 .812629307e+09                   4
BIN25AJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98303999
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869678823e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987939310e+11 .812629307e+09                   4
BIN25AJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     98303999
 .485549182e+09 .776062114e+06-.286822983e+03 .477740005e-01-.297195711e-05    2
-.869678823e+11-.250206781e+10-.140855400e+09 .213985655e+07-.675692266e+03    3
-.790697240e+00 .486960330e-03 .987939310e+11 .812629307e+09                   4
BIN25BJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65535999
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985634e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016860e+11 .726140704e+09                   4
BIN25BJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65535999
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985634e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016860e+11 .726140704e+09                   4
BIN25BJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     65535999
 .458257901e+09 .732441964e+06-.270701515e+03 .450887658e-01-.280491225e-05    2
-.138985634e+12-.243024799e+10-.137907599e+09 .200703096e+07-.540292703e+03    3
-.864558013e+00 .497990623e-03 .370016860e+11 .726140704e+09                   4
BIN25CJaggI             C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384000
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012262e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556866802e+11 .596407805e+09                   4
BIN25CJaggII            C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384000
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012262e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556866802e+11 .596407805e+09                   4
BIN25CJaggIII           C   0H   0          G   300.00   4000.00  1000.00      1&
C    327680000 H     16384000
 .417320981e+09 .667011741e+06-.246519312e+03 .410609140e-01-.255434495e-05    2
-.217012262e+12-.232251827e+10-.133485899e+09 .180779258e+07-.337193359e+03    3
-.975349173e+00 .514536064e-03-.556866802e+11 .596407805e+09                   4
END
