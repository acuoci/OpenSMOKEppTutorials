! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: TOT2003.THERM
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 3/24/2020

THERMO ALL
270.   1000.   3500. 
AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013931e+00-3.98290200e-07 3.45886082e-10-1.18293971e-13 1.38553174e-17    2
-7.45407891e+02 4.37897362e+00 2.49974489e+00 1.52569132e-06-3.17359231e-09    3
 2.74307057e-12-8.58511922e-16-7.45343207e+02 4.38079817e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811579e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324662e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42576298e-07 4.63926302e-10-1.57302170e-13 1.82971406e-17    2
-7.45426807e+02 9.27648988e-01 2.49964853e+00 2.08151569e-06-4.16682427e-09    3
 3.47465907e-12-1.04992675e-15-7.45332012e+02 9.30248556e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873259e-03 1.24226233e-06-4.19011898e-10 4.75543793e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529274e-03-1.27163634e-05    3
 1.28749173e-08-4.70027749e-12-9.43236614e+02-5.12231102e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406828e-07 6.39345346e-10-2.12551791e-13 2.44479191e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164046e-06-5.92759759e-09    3
 4.87810165e-12-1.45539320e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556201e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740147e-03 9.80122558e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959644e-04 1.33918546e-07-3.85875896e-11 4.38918689e-15    2
 2.92061519e+04 4.48358519e+00 3.14799201e+00-3.11174065e-03 6.18137897e-06    3
-5.63808798e-09 1.94866016e-12 2.91309118e+04 2.13446549e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218862e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710799e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805705e-03 5.06678941e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255381e+00 1.87486886e-03-8.59711926e-07 1.91200070e-10-1.67855286e-14    2
-1.41723335e+04 7.41443560e+00 3.75723891e+00-2.14465241e-03 5.42079005e-06    3
-4.17025963e-09 1.11901127e-12-1.43575530e+04 2.79976799e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876468e+00 2.62914704e-03-9.30606462e-07 1.43892920e-10-7.62581414e-15    2
-4.90562639e+04-2.34976452e+00 2.31684347e+00 9.22755036e-03-7.75654093e-06    3
 3.28225360e-09-5.48722482e-13-4.83626067e+04 1.00786234e+01                   4
HOCO                    H   1C   1O   2     G    200.00   3500.00 1570.00      1
 5.88810541e+00 3.28985507e-03-9.88703861e-07 1.12295277e-10-2.32818718e-15    2
-2.40914384e+04-5.05613727e+00 2.36661498e+00 1.22618052e-02-9.56063074e-06    3
 3.75217930e-09-5.81927554e-13-2.29856904e+04 1.35214769e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346405e-01 1.23697845e-02-4.99807922e-06 1.04392765e-09-8.62897416e-14    2
-9.58982501e+03 1.61752775e+01 5.23967335e+00-1.46835123e-02 5.29732711e-05    3
-5.41668822e-08 1.96318566e-11-1.02526308e+04-4.97649748e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805104e+00 6.15233477e-03-2.21179349e-06 3.74402648e-10-2.48151349e-14    2
 1.65862829e+04 5.77899818e+00 3.47829310e+00 3.54764773e-03 1.47408440e-06    3
-1.94375955e-09 5.21921232e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272972e+00 3.55431388e-03-1.28768523e-06 2.21273744e-10-1.48738147e-14    2
 4.62073492e+04 6.64284652e+00 3.76489460e+00 1.43839191e-03 4.75583077e-07    3
-4.31788591e-10 7.58292874e-14 4.58645699e+04 1.48953153e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468307e-03-1.35589914e-06 2.74980411e-10-2.36795472e-14    2
 5.06429079e+04 6.11646383e+00 4.18185434e+00-2.21134314e-03 7.71527541e-06    3
-5.95950381e-09 1.58314628e-12 5.03669407e+04-7.03002602e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472531e+00 3.92839476e-05-6.70014980e-08 3.71818694e-11-5.07306885e-15    2
 8.54504422e+04 4.79314254e+00 2.54495192e+00-2.47725281e-04 5.48018277e-07    3
-5.48551250e-10 2.04117331e-13 8.54434105e+04 4.56874273e+00                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990128e+00 2.16985238e-03-7.07637885e-07 1.23973494e-10-9.56348515e-15    2
 7.11059412e+04 8.77326061e+00 3.77264332e+00-1.58547350e-03 2.83512238e-06    3
-1.36146058e-09 2.23995332e-13 7.06312492e+04 8.79407904e-01                   4
CH3O2H                  C   1H   4O   2     G    300.00   3500.00 1090.00      1
 7.33435519e+00 9.33238534e-03-3.40995713e-06 5.79327692e-10-3.79241109e-14    2
-1.81046374e+04-1.19553974e+01 7.70006797e-01 3.34217373e-02-3.65604414e-05    3
 2.08548532e-08-4.68827401e-12-1.66736094e+04 2.02794895e+01                   4
CH3O2                   C   1H   3O   2     G    300.00   3500.00 1800.00      1
 5.64141817e+00 8.74328281e-03-3.21961406e-06 5.43695218e-10-3.45015008e-14    2
-1.19010148e+03-3.41914683e+00 1.44289632e+00 1.80733314e-02-1.09946545e-05    3
 3.42333984e-09-4.34452142e-13 3.21366390e+02 1.93041293e+01                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701530e+00 1.21538353e-02-5.02107031e-06 1.01068070e-09-8.18460823e-14    2
-2.57693409e+04 9.47420540e+00 8.47330479e-01 1.63086904e-02-8.48344961e-06    3
 2.29304341e-09-2.59952013e-13-2.50962544e+04 1.95933297e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238062e+00 5.90227637e-03-1.80340720e-06 2.13335009e-10-5.61816409e-15    2
-7.86252225e+01-7.49173677e+00 8.89660985e-01 1.70119767e-02-1.13807351e-05    3
 3.88280928e-09-5.32841479e-13 1.60316121e+03 1.85001134e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534950e+00 6.02727059e-03-2.11386821e-06 3.36085905e-10-2.00987482e-14    2
-4.03584143e+03-1.57524073e+00 2.34821579e+00 1.39600168e-02-1.08632206e-05    3
 4.62498416e-09-8.08499162e-13-3.30222106e+03 1.22661977e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335652e+00 1.00905183e-02-5.12952562e-06 1.25425207e-09-1.19639109e-13    2
-1.39080170e+04 1.59916144e+01 4.32621296e+00-7.01151853e-03 3.15176961e-05    3
-3.36478638e-08 1.23454023e-11-1.43270169e+04 2.62028902e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278258e-03-2.69184211e-06 7.21357798e-10-7.43521409e-14    2
 4.05725330e+03 1.07450933e+01 4.03483979e+00-2.15836864e-03 1.18233875e-05    3
-1.18459406e-08 4.00593954e-12 3.83636392e+03 4.20008770e+00                   4
HO2CHO                  C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230825e+01 4.43559488e-03-1.56185338e-06 2.43413972e-10-1.38379570e-14    2
-3.81313380e+04-2.33591553e+01 2.47434345e+00 2.16898555e-02-1.63512196e-05    3
 5.87745825e-09-8.18701426e-13-3.54892793e+04 1.72835404e+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473661e+00 8.42765725e-03-3.84722250e-06 8.63389842e-10-7.73674422e-14    2
-4.73118221e+04 5.12933885e+00 1.85206266e+00 1.27447105e-02-7.44476686e-06    3
 2.19581368e-09-2.62426309e-13-4.66124595e+04 1.56434956e+01                   4
OCHO                    C   1O   2H   1     G    200.00   3500.00  700.00      1
 2.58373953e+00 8.99565940e-03-4.55939787e-06 1.11902584e-09-1.07899898e-13    2
-1.67164582e+04 1.34890938e+01 4.25809175e+00-5.72067562e-04 1.59428742e-05    3
-1.84069475e-08 6.86566202e-12-1.69508675e+04 6.00851172e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959141e+00 1.57445261e-02-5.96197393e-06 1.06867182e-09-7.61012340e-14    2
-1.25948053e+04-1.43089412e+00-2.41778724e-01 2.53475709e-02-1.39645112e-05    3
 4.03257452e-09-4.87754387e-13-1.10391121e+04 2.19572625e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791360e+00 1.11042800e-02-3.71281686e-06 5.47665571e-10-2.89412604e-14    2
 1.17176215e+04-4.91382513e+00 6.75421801e-01 2.11542617e-02-1.20878017e-05    3
 3.64951180e-09-4.59753237e-13 1.33457186e+04 1.95628439e+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   3500.00 1450.00      1
 1.00876750e+01 1.40221806e-02-4.79128015e-06 7.15474133e-10-3.78163629e-14    2
-2.40669299e+04-2.56733582e+01-5.77204918e-01 4.34425389e-02-3.52261336e-05    3
 1.47085102e-08-2.45040879e-12-2.09741147e+04 2.97412031e+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   3500.00 1480.00      1
 9.29919683e+00 1.29334624e-02-4.54028592e-06 7.01327861e-10-3.92078228e-14    2
-7.64002445e+03-2.14311736e+01 2.00183268e-01 3.75253910e-02-2.94645378e-05    3
 1.19284684e-08-1.93568426e-12-4.94671644e+03 2.60335034e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402718e+00 9.50595350e-03-3.15129261e-06 4.53052074e-10-2.23949159e-14    2
 3.97229102e+03-3.77420905e+00-6.02932450e-02 2.08133970e-02-1.34307867e-05    3
 4.60638301e-09-6.51687481e-13 5.51151676e+03 2.10642172e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728376e+00 7.47581588e-03-2.58984227e-06 4.05265795e-10-2.35022721e-14    2
 3.38403785e+04 1.51958751e+00 1.23421214e+00 1.56222204e-02-1.10171572e-05    3
 4.27989337e-09-6.91541509e-13 3.46967692e+04 1.68637048e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267454e+00 5.47212830e-03-2.03181542e-06 3.75019116e-10-2.77049062e-14    2
 2.58626597e+04-2.43835921e+00 7.70536907e-01 2.37107998e-02-3.66622044e-05    3
 2.95989761e-08-9.27579255e-12 2.64317975e+04 1.40907683e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788257e+00 4.21328989e-03-1.58936946e-06 2.68739191e-10-1.73346359e-14    2
 6.72874491e+04 5.32512367e+00 4.60873599e+00 1.42766785e-03 8.54158643e-07    3
-6.83903344e-10 1.21940589e-13 6.68801772e+04-1.05894068e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490827e+00 1.39762977e-02-4.67366748e-06 6.82063684e-10-3.47025038e-14    2
-3.18909574e+04-1.38313071e+01-4.22291411e-01 3.35894614e-02-2.32937596e-05    3
 8.53864266e-09-1.27783209e-12-2.94428423e+04 2.70882146e+01                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957255e+00 2.35453825e-02-1.23415273e-05 3.08911893e-09-2.98016648e-13    2
-3.10347953e+03 1.69410913e+01 3.27852943e+00 1.44656289e-02 7.11508755e-06    3
-1.54409905e-08 6.31987957e-12-3.32593350e+03 9.84203392e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479680e+00 1.17471700e-02-4.06239751e-06 6.31554725e-10-3.61645074e-14    2
-6.24418450e+03-9.60110092e+00 1.82077785e+00 2.63431399e-02-1.89562444e-05    3
 7.38613379e-09-1.18490244e-12-4.66716293e+03 1.83437446e+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1500.00      1
 6.63757422e+00 1.19924585e-02-4.07718738e-06 6.22004997e-10-3.47508084e-14    2
-9.66525354e+03-7.65007787e+00 1.23305393e+00 2.64045127e-02-1.84892415e-05    3
 7.02736239e-09-1.10231037e-12-8.04389745e+03 2.06149529e+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   3500.00 1440.00      1
 9.66417632e+00 1.29483231e-02-4.44318337e-06 6.83406482e-10-3.84804393e-14    2
 1.86599132e+03-2.38806241e+01 2.23212418e+00 3.35929124e-02-2.59479639e-05    3
 1.06393234e-08-1.76693824e-12 4.00642234e+03 1.46847781e+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   3500.00 1520.00      1
 6.04215804e+00 1.11433647e-02-3.80167462e-06 5.65226940e-10-2.94248186e-14    2
-9.44151524e+03-1.02352918e+01-2.19672856e+00 3.28246452e-02-2.51976751e-05    3
 9.94943769e-09-1.57288053e-12-6.93689371e+03 3.29622805e+01                   4
C2H3O1-2                C   2H   3O   1     G    200.00   3500.00 1800.00      1
 7.60993625e+00 6.11300596e-03-1.59366937e-06 1.28294159e-10 2.98968068e-15    2
 1.61313302e+04-1.70584528e+01 7.34197746e-02 2.28608204e-02-1.55501814e-05    3
 5.29737268e-09-7.14937891e-13 1.88444761e+04 2.37307466e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195371e+00 1.06589270e-02-3.75190329e-06 6.00731628e-10-3.66603824e-14    2
-2.30621355e+04-8.31408577e+00 9.75916637e-01 2.23167871e-02-1.34667868e-05    3
 4.19883662e-09-5.36397187e-13-2.11735621e+04 2.00785613e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 6.07689016e+00 8.12979339e-03-2.81854999e-06 4.38698307e-10-2.55171837e-14    2
-4.06801047e+03-6.15492453e+00 1.47388064e+00 1.83587034e-02-1.13426417e-05    3
 3.59576931e-09-4.63999267e-13-2.41092705e+03 1.87575232e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703792e+00 7.91358604e-03-2.83605891e-06 4.62112655e-10-2.83231297e-14    2
-1.16170812e+03-8.37157286e+00 7.37868281e-01 2.50454357e-02-2.20135026e-05    3
 1.00031294e-08-1.80836357e-12 3.76389339e+02 2.09962837e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523628e+00 6.46841658e-03-2.33588414e-06 3.83408110e-10-2.36897850e-14    2
-8.05944305e+03-4.61154403e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226119e-09-9.59140718e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420513e+00 3.89116779e-03-1.41168608e-06 2.35668533e-10-1.49424971e-14    2
 1.94026782e+04-4.94089647e+00 3.33028661e+00 1.20351629e-02-1.14247949e-05    3
 5.70731267e-09-1.13618105e-12 2.00087543e+04 7.53650387e+00                   4
HCOOH                   C   1H   2O   2     G    300.00   3500.00 1640.00      1
 5.21581644e+00 5.48253641e-03-1.72756111e-06 2.25438490e-10-8.81949912e-15    2
-4.56198641e+04-2.59494560e+00 1.19691275e+00 1.52847405e-02-1.06929917e-05    3
 3.86992247e-09-5.64381082e-13-4.43016637e+04 1.87820781e+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483420e-03 1.65900439e-06-8.55133989e-10 9.82287244e-14    2
-2.73756816e+04-4.36816973e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH2OHCHO                C   2H   4O   2     G    300.00   3500.00 1800.00      1
 8.91045186e+00 9.14305837e-03-2.53718677e-06 2.39203912e-10 8.50819938e-16    2
-4.09945450e+04-1.84179622e+01 1.56305396e+00 2.54706093e-02-1.61434792e-05    3
 5.27857147e-09-6.99061342e-13-3.83494818e+04 2.13476880e+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   3500.00 1570.00      1
 9.97760259e+00 4.26981223e-03-1.12729433e-06 7.37809055e-11 5.98360578e-15    2
-2.96900177e+04-2.75230973e+01 7.08345765e-01 2.78857532e-02-2.36902952e-05    3
 9.65467301e-09-1.51963616e-12-2.67794711e+04 2.13768445e+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319128e-02-1.90892866e-05    3
 5.92848299e-09-7.42884555e-13-1.63833552e+04 6.70139035e+00                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772145e-02-4.04888397e-06 6.94756696e-10-4.56573670e-14    2
-7.51809422e+04-3.74730276e+01-2.33886892e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164715e-12-7.15304886e+04 3.67067395e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 5.02910657e+00-2.87377519e-02 6.15808970e-05-2.98073518e-08 4.29774802e-12    2
-4.07046731e+04 1.82412181e+01 2.12034974e-07-1.31715123e-09 2.87530013e-12    3
 2.88411189e-08-1.66481344e-11-4.00005982e+04 4.07099930e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849390e-09-3.11411020e-13    2
-2.07588781e+04 1.60124236e+01 4.66126893e+00 9.68655552e-03 1.14715528e-05    3
-1.83003965e-08 7.03409940e-12-2.10634335e+04 6.60518516e+00                   4
C3H8                    C   3H   8          G    300.00   3500.00 1690.00      1
 8.33847007e+00 1.79340922e-02-5.80534981e-06 7.91037708e-10-3.43401227e-14    2
-1.70816233e+04-2.27461799e+01-1.38651266e+00 4.09518028e-02-2.62352705e-05    3
 8.85017800e-09-1.22652064e-12-1.37945792e+04 2.92742161e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1800.00      1
 6.05951251e+00 1.82035621e-02-6.54041321e-06 1.09272144e-09-7.13189353e-14    2
 7.29671818e+03-6.80793083e+00-6.08211221e-01 3.30207259e-02-1.88880497e-05    3
 5.66592015e-09-7.06485424e-13 9.69709872e+03 2.92791809e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1590.00      1
 7.21724982e+00 1.65877265e-02-5.58902439e-06 8.31338515e-10-4.40999325e-14    2
 8.50975633e+03-1.26938767e+01-1.37086178e-01 3.50892007e-02-2.30432453e-05    3
 8.14967015e-09-1.19478101e-12 1.08484352e+04 2.61969991e+01                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755201e+00 1.65820017e-02-6.59972302e-06 1.29512916e-09-1.03784375e-13    2
-3.79456071e+02-1.05616187e+01-8.55987188e-02 3.08112255e-02-1.84574096e-05    3
 5.68686491e-09-7.13747674e-13 1.92567819e+03 2.40935687e+01                   4
C3H5-A                  C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877792e+00 1.04611885e-02-3.15379708e-06 3.85306884e-10-1.26413689e-14    2
 1.71766363e+04-2.28181758e+01-3.57888096e-01 3.27028536e-02-2.40053580e-05    3
 9.07345729e-09-1.37016487e-12 2.00235695e+04 2.42845603e+01                   4
C3H5-S                  C   3H   5          G    300.00   3500.00 1800.00      1
 6.52599516e+00 1.37686655e-02-5.50691342e-06 1.07278366e-09-8.39560017e-14    2
 2.86430050e+04-9.99635700e+00 1.54227621e+00 2.48435965e-02-1.47360226e-05    3
 4.49097224e-09-5.58704416e-13 3.04371438e+04 1.69765696e+01                   4
C3H5-T                  C   3H   5          G    300.00   3500.00  770.00      1
 1.49331935e+00 2.33788729e-02-1.18550710e-05 2.86552470e-09-2.68203790e-13    2
 2.87117775e+04 1.76892214e+01 2.52238869e+00 1.80330581e-02-1.44114618e-06    3
-6.15086046e-09 2.65919399e-12 2.85533009e+04 1.29935191e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079978e+00 1.37589661e-02-5.15319199e-06 9.32421983e-10-6.74695911e-14    2
 7.77376170e+03-2.10036658e+01 9.27196847e-01 3.40908988e-02-2.40959865e-05    3
 8.77622923e-09-1.28545208e-12 1.04088818e+04 2.23747992e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1550.00      1
 9.00938222e+00 1.57632590e-02-5.29374355e-06 7.64253417e-10-3.74126438e-14    2
-1.56669515e+04-2.44960178e+01-1.88321638e+00 4.38731909e-02-3.24969034e-05    3
 1.24645372e-08-1.92455519e-12-1.22902459e+04 3.28282089e+01                   4
CH3CHCHO                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 6.70347362e+00 1.89922318e-02-9.18109977e-06 2.14445657e-09-1.96154637e-13    2
-6.21094363e+03-1.05801331e+01 2.92067498e-01 3.32398010e-02-2.10540741e-05    3
 6.54185446e-09-8.06904344e-13-3.90283743e+03 2.41197343e+01                   4
AC4H7OOH                C   4H   8O   2     G    300.00   3500.00 1660.00      1
 1.22738272e+01 2.55483383e-02-9.81265077e-06 1.82078670e-09-1.35039880e-13    2
-1.24525960e+04-3.36837474e+01 1.60151447e+00 5.12647544e-02-3.30503762e-05    3
 1.11532065e-08-1.54052480e-12-8.90938817e+03 2.32129081e+01                   4
CH3CHCO                 C   3H   4O   1     G    300.00   3500.00 1280.00      1
 6.99681463e+00 1.49445085e-02-6.71568578e-06 1.45955079e-09-1.25293200e-13    2
-1.29366480e+04-1.07908059e+01 1.50068777e+00 3.21199049e-02-2.68431035e-05    3
 1.19425808e-08-2.17276001e-12-1.15296395e+04 1.70816035e+01                   4
AC3H5OOH                C   3H   6O   2     G    298.00   3500.00 1800.00      1
 1.36957657e+01 1.27112963e-02-4.21186263e-06 6.49030109e-10-3.94931202e-14    2
-1.11479407e+04-4.31791016e+01 4.22354618e+00 3.37606729e-02-2.17530098e-05    3
 7.14575129e-09-9.41815506e-13-7.73794171e+03 8.08652616e+00                   4
C3H6OH1-2               C   3H   7O   1     G    300.00   3500.00 1800.00      1
 8.46016352e+00 1.89669003e-02-7.38013554e-06 1.39189577e-09-1.05413394e-13    2
-1.21581707e+04-1.51603324e+01 4.08605477e-01 3.68592515e-02-2.22904282e-05    3
 6.91422639e-09-8.72403758e-13-9.25960980e+03 2.84163793e+01                   4
C3H6OH2-1               C   3H   7O   1     G    300.00   3500.00 1590.00      1
 8.99548234e+00 1.75103792e-02-6.94615357e-06 1.37004323e-09-1.07539337e-13    2
-1.65436320e+04-1.93287236e+01 1.31207693e+00 3.68397010e-02-2.51813628e-05    3
 9.01583327e-09-1.30970758e-12-1.41003090e+04 2.13023225e+01                   4
HOC3H6O2                C   3H   7O   3     G    300.00   3500.00 1480.00      1
 1.24409055e+01 2.15172909e-02-8.97737594e-06 1.82414691e-09-1.48047122e-13    2
-3.10315628e+04-3.23089026e+01 2.93449048e+00 4.72103044e-02-3.50175923e-05    3
 1.35539741e-08-2.12943685e-12-2.82176640e+04 1.72809693e+01                   4
SC3H5OH                 C   3H   6O   1     G    300.00   3500.00 1260.00      1
 7.83167544e+00 1.85990426e-02-7.98421836e-06 1.67672190e-09-1.40411942e-13    2
-2.22362405e+04-1.56369776e+01-5.71229678e-02 4.36428470e-02-3.77982713e-05    3
 1.74513531e-08-3.27029908e-12-2.02482633e+04 2.42451084e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00 1630.00      1
 9.39463114e+00 1.51343106e-02-4.86246276e-06 6.64177249e-10-2.94552530e-14    2
-2.20582199e+04-2.45922026e+01 4.73537667e-01 3.70265645e-02-2.50087087e-05    3
 8.90395064e-09-1.29322418e-12-1.91499434e+04 2.28055845e+01                   4
CH2CCH2OH               C   3H   5O   1     G    300.00   3500.00 1800.00      1
 7.15397365e+00 1.62590933e-02-7.06959971e-06 1.52062107e-09-1.30983749e-13    2
 1.01359982e+04-8.36739478e+00 2.39300609e+00 2.68390212e-02-1.58862063e-05    3
 4.78603091e-09-5.84512894e-13 1.18499465e+04 1.73999548e+01                   4
C3H4-P                  C   3H   4          G    300.00   3500.00 1570.00      1
 6.45797858e+00 1.06371316e-02-3.61161722e-06 5.39412691e-10-2.85851275e-14    2
 1.94136786e+04-1.10770989e+01 1.72714322e+00 2.26902153e-02-1.51273023e-05    3
 5.42930020e-09-8.07229635e-13 2.08991609e+04 1.38804115e+01                   4
C3H4-A                  C   3H   4          G    300.00   3500.00 1420.00      1
 6.37608366e+00 1.10282079e-02-3.89476312e-06 6.16686076e-10-3.59564768e-14    2
 2.00917847e+04-1.13283006e+01 5.08248696e-01 2.75573205e-02-2.13550933e-05    3
 8.81402419e-09-1.47914981e-12 2.17582498e+04 1.90382079e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057762e+00 1.05635747e-02-4.84060952e-06 1.09040068e-09-9.80036130e-14    2
 4.00565408e+04-5.04125059e+00 1.75584147e+00 2.95861278e-02-3.88094543e-05    3
 2.80498013e-08-8.12163476e-12 4.07276565e+04 1.35345464e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00 1260.00      1
 6.42043189e+00 6.05128866e-03-2.30888141e-06 4.10631875e-10-2.84293474e-14    2
 6.08598164e+04-8.32404334e+00 2.15397882e+00 1.95955841e-02-1.84330427e-05    3
 8.94193413e-09-1.72114805e-12 6.19349626e+04 1.32451538e+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1710.00      1
 9.33264604e+00 1.46861072e-02-4.56011955e-06 5.69518135e-10-1.90908109e-14    2
-2.69164882e+04-2.52385565e+01-9.86882752e-02 3.67477080e-02-2.39124009e-05    3
 8.11426720e-09-1.12212430e-12-2.36909719e+04 2.53220280e+01                   4
CH2CH2CHO               C   3H   5O   1     G    300.00   3500.00  700.00      1
 1.38640400e+00 2.84363938e-02-1.56688640e-05 4.07196321e-09-4.03232083e-13    2
 6.14151634e+02 2.19844218e+01 2.41071832e+00 2.25831692e-02-3.12623980e-06    3
-7.87339320e-09 3.86296664e-12 4.70747631e+02 1.74080446e+01                   4
RALD3                   C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180078e-02-2.61696720e-05 6.65382129e-09-6.35305357e-13    2
-2.14966001e+03 5.90959840e+01 7.04072886e+00-2.01204450e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381685e+00                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597839e+00 1.12038372e-02-3.67974365e-06 5.08180252e-10-2.25803375e-14    2
-1.23719484e+04-2.08137560e+01 8.18908043e-01 3.22215131e-02-2.33838148e-05    3
 8.71820989e-09-1.30539747e-12-9.68168587e+03 2.36968522e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00 1790.00      1
 9.79507855e+00 1.35932465e-02-4.01642284e-06 4.43034305e-10-7.94380246e-15    2
-3.07542949e+04-2.70699391e+01-7.54581368e-03 3.54985524e-02-2.23728244e-05    3
 7.27968292e-09-9.62782995e-13-2.72449554e+04 2.59292980e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1590.00      1
 8.40473847e+00 1.29432044e-02-4.25667366e-06 6.02254911e-10-2.86748418e-14    2
-7.89528923e+03-1.63899805e+01 1.00367440e+00 3.15622335e-02-2.18217955e-05    3
 7.96708586e-09-1.18666713e-12-5.54175085e+03 2.27480006e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14851999e-06-5.94424210e-11 5.32964638e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
PC4H9                   C   4H   9          G    300.00   3500.00  950.00      1
 3.94763006e+00 3.16286394e-02-1.12984867e-05 1.11637450e-09 5.54031605e-14    2
 6.05554723e+03 7.76350061e+00-2.76188385e-01 4.94131381e-02-3.93792741e-05    3
 2.08221903e-08-5.13033783e-12 6.85807273e+03 2.79243295e+01                   4
SC4H9                   C   4H   9          G    300.00   3500.00  850.00      1
 3.40122928e+00 3.20901863e-02-1.12255470e-05 9.71712110e-10 8.30726274e-14    2
 4.66283101e+03 1.05291639e+01 2.36336421e-01 4.69837998e-02-3.75083943e-05    3
 2.15857099e-08-5.97986791e-12 5.20086280e+03 2.52835874e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955795e+00 3.23747266e-02-1.18655436e-05 1.37455177e-09 1.57073481e-14    2
-1.97025810e+04-6.34483426e+00-1.85965329e+00 5.58007941e-02-3.97537191e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H9                   C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221490e-06 8.09648920e-10 4.02033223e-14    2
 3.37759297e+03-1.61084037e+01-1.15582377e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
TC4H9                   C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871689e+00 2.55264450e-02-8.65284049e-06 8.24419700e-10 3.80550657e-14    2
 8.35470579e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397361e-05    3
 1.42467509e-08-2.35878980e-12 3.41363196e+03 3.01901373e+01                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385767e+03-1.72949366e+01 7.17301599e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035733e-13-3.72372397e+03 2.01415164e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177117e+00 3.67769037e-02-1.77031337e-05 3.74786266e-09-2.92191284e-13    2
 1.31214242e+04 2.00120540e+01 3.86130010e+00 2.14653098e-02 1.51074247e-05    3
-2.75002882e-08 1.08678626e-11 1.27462902e+04 8.04059663e+00                   4
IC4H7O                  C   4H   7O   1     G    300.00   3500.00 1800.00      1
 1.18822163e+01 1.89918532e-02-7.42296498e-06 1.41442848e-09-1.08683660e-13    2
 1.15971319e+03-3.56333819e+01 1.50010972e+00 4.20632012e-02-2.66490883e-05    3
 8.53521488e-09-1.09768177e-12 4.89727156e+03 2.05567447e+01                   4
C4H8-1                  C   4H   8          G    300.00   3500.00 1800.00      1
 1.03330449e+01 1.99470428e-02-7.40538998e-06 1.30472507e-09-9.09598189e-14    2
-5.56551437e+03-3.07722296e+01-6.91489888e-01 4.44460090e-02-2.78211951e-05    3
 8.86613439e-09-1.14115556e-12-1.59668184e+03 2.88948525e+01                   4
C4H8-2                  C   4H   8          G    300.00   3500.00 1800.00      1
 5.15907399e+00 2.89997694e-02-1.32974598e-05 2.96139017e-09-2.60424474e-13    2
-4.76704683e+03-3.39008062e+00 5.60608454e-01 3.92185817e-02-2.18131368e-05    3
 6.11534459e-09-6.98473698e-13-3.11159924e+03 2.14977742e+01                   4
C4H71-3                 C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017754e+00 1.98466503e-02-6.37614061e-06 5.28652768e-10 3.81103734e-14    2
 1.19533850e+04-1.83767119e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
C4H71-4                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075605e-06 3.82147970e-10 5.73994809e-14    2
 1.98988324e+04-1.80212793e+01-3.29329052e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
C4H71-O                 C   4H   7O   1     G    300.00   3500.00 1600.00      1
 1.37371777e+01 1.70982846e-02-6.55972544e-06 1.21466090e-09-8.98269615e-14    2
-3.28789072e+01-4.64105970e+01-1.48200925e+00 5.51462520e-02-4.22296948e-05    3
 1.60771481e-08-2.41209059e-12 4.83726091e+03 3.41662556e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872521e+00 1.50139591e-02-5.06688177e-06 7.84148097e-10-4.70262839e-14    2
 8.60829987e+03-2.47389586e+01 4.65225109e-01 3.46661815e-02-2.14437338e-05    3
 6.84964885e-09-8.89456944e-13 1.17919599e+04 2.31239087e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794386e-03 4.88814514e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742308e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777119e+00 1.26498258e-02-4.62248950e-06 7.81217082e-10-5.07629107e-14    2
 3.13366016e+04-1.49692661e+01 7.13119716e-01 3.41836288e-02-2.96617954e-05    3
 1.37214268e-08-2.55855550e-12 3.31283217e+04 2.03030643e+01                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590364e-03 1.80568200e-06-9.30237204e-10 1.18077198e-13    2
 6.01811751e+04-4.25791500e+01 2.34662666e+00 2.83894138e-02-2.35278181e-05    3
 9.69177543e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00  720.00      1
 7.13414735e+00 1.00526308e-02-4.84819206e-06 1.14884604e-09-1.07722834e-13    2
 5.27577824e+04-1.36443516e+01-4.34754087e-01 5.21020832e-02-9.24512179e-05    3
 8.22627589e-08-2.82722759e-11 5.38477042e+04 2.03848077e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055544e+01 1.99961045e-02-7.07935460e-06 1.10673028e-09-6.24178899e-14    2
 4.11452290e+03-4.24445091e+01-6.99882110e+00 7.24907868e-02-6.29247613e-05    3
 2.75111779e-08-4.74405754e-12 9.33275680e+03 5.31863191e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152220e+01 1.47750067e-02-3.90939181e-06 2.82308156e-10 1.62511622e-14    2
 1.91167581e+04-5.54965184e+01-3.67012639e+00 6.11476948e-02-4.84985149e-05    3
 1.93374890e-08-3.03746371e-12 2.47593868e+04 3.97971310e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331261e+01 1.77269649e-02-6.33615682e-06 1.00236865e-09-5.75481750e-14    2
 3.49856300e+04-3.80075865e+01-6.76261385e+00 6.95132669e-02-6.22206553e-05    3
 2.78054854e-08-4.87825263e-12 3.99884457e+04 5.47375207e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786764e+01 1.28174257e-02-3.11961936e-06 1.29368393e-10 2.76958521e-14    2
 9.43770579e+03-5.26289052e+01-4.05866643e+00 5.60992486e-02-4.29495178e-05    3
 1.64197154e-08-2.47082363e-12 1.51874796e+04 4.10783319e+01                   4
C5H5                    C   5H   5          G    300.00   3500.00  700.00      1
 4.01652588e+00 2.68451887e-02-1.26423015e-05 2.78092323e-09-2.35299425e-13    2
 2.91110159e+04 1.44025731e+00-2.58737467e+00 6.45817633e-02-9.35063898e-05    3
 7.97943407e-08-2.77400914e-11 3.00355619e+04 3.09448142e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1470.00      1
 1.21408016e+01 2.34281374e-02-7.98702759e-06 1.18908391e-09-6.20202054e-14    2
 7.23040214e+03-4.21606537e+01-5.49894699e+00 7.14274534e-02-5.69659215e-05    3
 2.34017342e-08-3.83968182e-12 1.24164882e+04 4.97368686e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248658e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987877e+01                   4
END
