!***********************************************************************
!SURFACE MECHANISM OF CH4 REFORMING AND OXIDATION OVER NI              *
!***********************************************************************
!****                                                                  *
!****     CH4 ON Ni - SURFACE MECHANISM                                *
!****
!****     Version 1.2  (March 2006)
!****
!****     V. Janardhanan, O. Deutschmann
!****     ITCP, University of Karlsruhe, Germany
!****     Contact: mail@detchem.com (O. Deutschmann)
!****
!****     NOTE: The mechanism Ni2005: E. Hecht, G.K. Gupta, H. Zhu. 
!****           A.M. Dean, R.J. Kee, L. Maier, O. Deutschmann.         *                    
!****           Applied Catalysis A: General 295 (2005) 40–51          
!****           adjusted for temperature range 500-2000°C for SOFC 
!****           applications
!****     Referenc:
!****     V.M. Janardhanan, O. Deutschmann. 
!****         Journal of Power Sources 162 (2006), 1192-1202
!****     www.detchem.com/mechanisms
!****
!****     Kinetic data:
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea
!****                                       (cm,mol,s)    -      J/mol
!****
!****
!****     Surface site density: 2.66E-9 mol/cm**2
!****
!****
!****     (SURFACE CHEMKIN format)
!****
!***********************************************************************

THERMO
   300.000  1000.000  3000.000

H2                121286H   2               G   300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633828E-06-0.09231578E-10 0.15827519E-14    2
-0.08350340E+04-0.13551101E+01 0.03298124E+02 0.08249441E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.10125209E+04-0.03294094E+02                   4
CH4           (adjust)  C   1H   4    0    0G   300.00   5000.00  1000.00      1
 1.68347883E+00 1.02372356E-02-3.87512864E-06 6.78558487E-10-4.50342312E-14    2
-1.00807871E+04 9.62339497E+00 7.78741479E-01 1.74766835E-02-2.78340904E-05    3
 3.04970804E-08-1.22393068E-11-9.82522852E+03 1.37221947E+01                   4
H2            (adjust)  H   2    0    0    0G   300.00   5000.00  1000.00      1
 3.06670950E+00 5.74737550E-04 1.39383190E-08-2.54835180E-11 2.90985740E-15    2
-8.65474120E+02-1.77984240E+00 3.35535140E+00 5.01361440E-04-2.30069080E-07    3
-4.79053240E-10 4.85225850E-13-1.01916260E+03-3.54772280E+00                   4
H2O           (adjust)  H   2O   1    0    0G   300.00   5000.00  1000.00      1
 2.61104720E+00 3.15631300E-03-9.29854380E-07 1.33315380E-10-7.46893510E-15    2
-2.98681670E+04 7.20912680E+00 4.16772340E+00-1.81149700E-03 5.94712880E-06    3
-4.86920210E-09 1.52919910E-12-3.02899690E+04-7.31354740E-01                   4
CO            (adjust)  C   1O   1    0    0G   300.00   5000.00  1000.00      1
 3.02507806E+00 1.44268852E-03-5.63082779E-07 1.01858133E-10-6.91095156E-15    2
-1.42683496E+04 6.10821772E+00 3.26245165E+00 1.51194085E-03-3.88175522E-06    3
 5.58194424E-09-2.47495123E-12-1.43105391E+04 4.84889698E+00                   4
CO2           (adjust)  C   1O   2    0    0G   300.00   5000.00  1000.00      1
 4.45362282E+00 3.14016873E-03-1.27841054E-06 2.39399667E-10-1.66903319E-14    2
-4.89669609E+04-9.55395877E-01 2.27572465E+00 9.92207229E-03-1.04091132E-05    3
 6.86668678E-09-2.11728009E-12-4.83731406E+04 1.01884880E+01                   4
O2            (adjust)  O   2    0    0    0G   300.00   5000.00  1000.00      1
 3.61221390E+00 7.48531660E-04-1.98206470E-07 3.37490080E-11-2.39073740E-15    2
-1.19781510E+03 3.67033070E+00 3.78371350E+00-3.02336340E-03 9.94927510E-06    3
-9.81891010E-09 3.30318250E-12-1.06381070E+03 3.64163450E+00                   4
AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2            (adjust)  N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
NI(s)         (adjust)  NI  1    0    0    0     300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O(s)        (adjust)  H   2O   1NI  1    0     500.00   2000.00 2000.00      1
 3.50421382E+00 6.68594839E-04 1.76268743E-06-1.17030152E-09 2.26185355E-13    2
-3.79129166E+04-1.05582534E+01 3.50421382E+00 6.68594839E-04 1.76268743E-06    3
-1.17030152E-09 2.26185355E-13-3.79129166E+04-1.05582534E+01                   4
H(s)          (adjust)  H   1NI  1    0    0     500.00   2000.00 2000.00      1
 1.38522354E+00-3.60291509E-05 1.01482878E-06-6.39234047E-10 1.26064639E-13    2
-5.45886573E+03-5.04262898E+00 1.38522354E+00-3.60291509E-05 1.01482878E-06    3
-6.39234047E-10 1.26064639E-13-5.45886573E+03-5.04262898E+00                   4
OH(s)         (adjust)  H   1O   1NI  1    0     500.00   2000.00 2000.00      1
 2.08905501E+00 1.71443903E-03-4.27838552E-07 9.11211411E-12 1.13760370E-14    2
-2.67334298E+04-3.86138841E+00 2.08905501E+00 1.71443903E-03-4.27838552E-07    3
 9.11211411E-12 1.13760370E-14-2.67334298E+04-3.86138841E+00                   4
CO(s)         (adjust)  C   1O   1NI  1    0     500.00   2000.00 2000.00      1
 1.04958397E+00 5.37825549E-03-3.51895909E-06 1.06323431E-09-1.12689240E-13    2
-2.73744388E+04 7.60559022E+00 1.04958397E+00 5.37825549E-03-3.51895909E-06    3
 1.06323431E-09-1.12689240E-13-2.73744388E+04 7.60559022E+00                   4
C(s)          (adjust)  C   1NI  1    0    0     500.00   2000.00 2000.00      1
-3.49330914E+00 5.23524687E-03-3.03308918E-06 6.55611035E-10-1.40966550E-14    2
-2.23124726E+03 7.68421239E+00-3.49330914E+00 5.23524687E-03-3.03308918E-06    3
 6.55611035E-10-1.40966550E-14-2.23124726E+03 7.68421239E+00                   4
CH3(s)        (adjust)  C   1H   3NI  1    0     500.00   2000.00 2000.00      1
-6.10760599E-01 8.61612510E-03-2.17714930E-06-6.63815294E-10 3.13819319E-13    2
-8.89792082E+03-2.00828704E+00-6.10760599E-01 8.61612510E-03-2.17714930E-06    3
-6.63815294E-10 3.13819319E-13-8.89792082E+03-2.00828704E+00                   4
CH2(s)        (adjust)  C   1H   2NI  1    0     500.00   2000.00 2000.00      1
-1.56917589E+00 7.30948876E-03-2.33683999E-06-2.63575385E-10 2.08877321E-13    2
 1.94307500E+03 4.44265982E+00-1.56917589E+00 7.30948876E-03-2.33683999E-06    3
-2.63575385E-10 2.08877321E-13 1.94307500E+03 4.44265982E+00                   4
CH(s)         (adjust)  C   1H   1NI  1    0     500.00   2000.00 2000.00      1
-2.52762352E+00 6.00297402E-03-2.49669461E-06 1.36758705E-10 1.03915796E-13    2
 9.56681068E+03 7.44010148E+00-2.52762352E+00 6.00297402E-03-2.49669461E-06    3
 1.36758705E-10 1.03915796E-13 9.56681068E+03 7.44010148E+00                   4
CH4(s)        (adjust)  C   1H   4NI  1    0     500.00   2000.00 2000.00      1
 3.47651462E-01 9.92277358E-03-2.01747493E-06-1.06404583E-09 4.18759375E-13    2
-1.38997273E+04-4.61646253E+00 3.47651462E-01 9.92277358E-03-2.01747493E-06    3
-1.06404583E-09 4.18759375E-13-1.38997273E+04-4.61646253E+00                   4
O(s)          (adjust)  O   1NI  1    0    0     500.00   2000.00 2000.00      1
 9.33885773E-01 1.49287485E-03-1.51153811E-06 7.60133452E-10-1.42499395E-13    2
-2.88011883E+04-3.47247502E+00 9.33885773E-01 1.49287485E-03-1.51153811E-06    3
 7.60133452E-10-1.42499395E-13-2.88011883E+04-3.47247502E+00                   4
CO2(s)        (adjust)  C   1O   2NI  1    0     500.00   2000.00 2000.00      1
 2.15782085E+00 8.85798101E-03-7.33295570E-06 3.01455469E-09-4.83617407E-13    2
-5.17211366E+04-3.96778204E-01 2.15782085E+00 8.85798101E-03-7.33295570E-06    3
 3.01455469E-09-4.83617407E-13-5.17211366E+04-3.96778204E-01                   4
HCO(s)        (adjust)  C   1H   1O   1NI  1     500.00   2000.00 2000.00      1
 1.42054865E+00 6.41898600E-03-3.25611216E-06 6.60406470E-10-1.25958802E-14    2
-1.72299589E+04-1.34060408E+00 1.42054865E+00 6.41898600E-03-3.25611216E-06    3
 6.60406470E-10-1.25958802E-14-1.72299589E+04-1.34060408E+00                   4

END
