! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: TOT2003.THERM
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 3/24/2020

THERMO ALL
270.   1000.   3500. 
AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013931e+00-3.98290200e-07 3.45886082e-10-1.18293971e-13 1.38553174e-17    2
-7.45407891e+02 4.37897362e+00 2.49974489e+00 1.52569132e-06-3.17359231e-09    3
 2.74307057e-12-8.58511922e-16-7.45343207e+02 4.38079817e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811579e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324662e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42576298e-07 4.63926302e-10-1.57302170e-13 1.82971406e-17    2
-7.45426807e+02 9.27648988e-01 2.49964853e+00 2.08151569e-06-4.16682427e-09    3
 3.47465907e-12-1.04992675e-15-7.45332012e+02 9.30248556e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873259e-03 1.24226233e-06-4.19011898e-10 4.75543793e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529274e-03-1.27163634e-05    3
 1.28749173e-08-4.70027749e-12-9.43236614e+02-5.12231102e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406828e-07 6.39345346e-10-2.12551791e-13 2.44479191e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164046e-06-5.92759759e-09    3
 4.87810165e-12-1.45539320e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556201e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740147e-03 9.80122558e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132646e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959644e-04 1.33918546e-07-3.85875896e-11 4.38918689e-15    2
 2.92061519e+04 4.48358519e+00 3.14799201e+00-3.11174065e-03 6.18137897e-06    3
-5.63808798e-09 1.94866016e-12 2.91309118e+04 2.13446549e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218862e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710799e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805705e-03 5.06678941e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
END
