! Examination of a Soot Model in Premixed Laminar Flames at Fuel-rich Conditions
! W. Pejpichestakul, E. Ranzi, M. Pelucchi, A. Frassoldati, A. Cuoci, A. Parente, T. Faravelli
! Proc. Combust. Inst. 37, 2019

THERMO ALL
270.   1000.   3500. 
AR                      AR  1               G    200.00   3500.00  820.00      1
 2.50013931e+00-3.98290225e-07 3.45886104e-10-1.18293978e-13 1.38553183e-17    2
-7.45407891e+02 4.37897362e+00 2.49974489e+00 1.52569140e-06-3.17359247e-09    3
 2.74307072e-12-8.58511967e-16-7.45343207e+02 4.38079817e+00                   4
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811580e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324661e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
HE                      HE  1               G    200.00   3500.00  850.00      1
 2.50020615e+00-5.42576318e-07 4.63926320e-10-1.57302176e-13 1.82971413e-17    2
-7.45426807e+02 9.27648988e-01 2.49964853e+00 2.08151575e-06-4.16682439e-09    3
 3.47465916e-12-1.04992678e-15-7.45332012e+02 9.30248556e-01                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873260e-03 1.24226233e-06-4.19011899e-10 4.75543794e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529275e-03-1.27163634e-05    3
 1.28749174e-08-4.70027750e-12-9.43236613e+02-5.12231094e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406872e-07 6.39345384e-10-2.12551804e-13 2.44479207e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164057e-06-5.92759783e-09    3
 4.87810185e-12-1.45539326e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556202e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740148e-03 9.80122560e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132645e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959648e-04 1.33918549e-07-3.85875908e-11 4.38918703e-15    2
 2.92061519e+04 4.48358518e+00 3.14799201e+00-3.11174063e-03 6.18137893e-06    3
-5.63808794e-09 1.94866014e-12 2.91309118e+04 2.13446550e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218863e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710800e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805704e-03 5.06678942e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255381e+00 1.87486886e-03-8.59711925e-07 1.91200070e-10-1.67855286e-14    2
-1.41723335e+04 7.41443560e+00 3.75723891e+00-2.14465241e-03 5.42079004e-06    3
-4.17025963e-09 1.11901127e-12-1.43575530e+04 2.79976799e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876468e+00 2.62914704e-03-9.30606462e-07 1.43892920e-10-7.62581413e-15    2
-4.90562639e+04-2.34976452e+00 2.31684347e+00 9.22755036e-03-7.75654093e-06    3
 3.28225360e-09-5.48722482e-13-4.83626067e+04 1.00786234e+01                   4
HOCO                    H   1C   1O   2     G    200.00   3500.00 1570.00      1
 5.88810541e+00 3.28985507e-03-9.88703861e-07 1.12295277e-10-2.32818717e-15    2
-2.40914384e+04-5.05613727e+00 2.36661498e+00 1.22618052e-02-9.56063074e-06    3
 3.75217930e-09-5.81927554e-13-2.29856904e+04 1.35214769e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346456e-01 1.23697844e-02-4.99807911e-06 1.04392761e-09-8.62897368e-14    2
-9.58982503e+03 1.61752773e+01 5.23967310e+00-1.46835107e-02 5.29732676e-05    3
-5.41668788e-08 1.96318554e-11-1.02526308e+04-4.97649641e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805104e+00 6.15233477e-03-2.21179349e-06 3.74402648e-10-2.48151348e-14    2
 1.65862829e+04 5.77899817e+00 3.47829310e+00 3.54764774e-03 1.47408439e-06    3
-1.94375954e-09 5.21921230e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272972e+00 3.55431388e-03-1.28768523e-06 2.21273744e-10-1.48738147e-14    2
 4.62073492e+04 6.64284652e+00 3.76489460e+00 1.43839191e-03 4.75583077e-07    3
-4.31788591e-10 7.58292874e-14 4.58645699e+04 1.48953153e+00                   4
CH2(S)                  C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468306e-03-1.35589913e-06 2.74980408e-10-2.36795469e-14    2
 5.06429079e+04 6.11646381e+00 4.18185434e+00-2.21134312e-03 7.71527537e-06    3
-5.95950378e-09 1.58314628e-12 5.03669407e+04-7.03002582e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472531e+00 3.92839476e-05-6.70014980e-08 3.71818694e-11-5.07306885e-15    2
 8.54504422e+04 4.79314254e+00 2.54495192e+00-2.47725281e-04 5.48018277e-07    3
-5.48551250e-10 2.04117331e-13 8.54434105e+04 4.56874273e+00                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990128e+00 2.16985238e-03-7.07637884e-07 1.23973494e-10-9.56348511e-15    2
 7.11059412e+04 8.77326061e+00 3.77264332e+00-1.58547350e-03 2.83512238e-06    3
-1.36146058e-09 2.23995331e-13 7.06312492e+04 8.79407904e-01                   4
CH3O2H                  C   1H   4O   2     G    300.00   3500.00 1090.00      1
 7.33435518e+00 9.33238537e-03-3.40995715e-06 5.79327700e-10-3.79241117e-14    2
-1.81046374e+04-1.19553973e+01 7.70006807e-01 3.34217372e-02-3.65604413e-05    3
 2.08548532e-08-4.68827399e-12-1.66736094e+04 2.02794894e+01                   4
CH3O2                   C   1H   3O   2     G    300.00   3500.00 1800.00      1
 5.64141817e+00 8.74328282e-03-3.21961407e-06 5.43695219e-10-3.45015008e-14    2
-1.19010148e+03-3.41914682e+00 1.44289632e+00 1.80733314e-02-1.09946545e-05    3
 3.42333984e-09-4.34452142e-13 3.21366390e+02 1.93041293e+01                   4
CH3OH                   C   1H   4O   1     G    300.00   3500.00 1800.00      1
 2.71701530e+00 1.21538353e-02-5.02107031e-06 1.01068070e-09-8.18460823e-14    2
-2.57693409e+04 9.47420541e+00 8.47330479e-01 1.63086904e-02-8.48344961e-06    3
 2.29304341e-09-2.59952013e-13-2.50962544e+04 1.95933297e+01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238062e+00 5.90227638e-03-1.80340720e-06 2.13335010e-10-5.61816419e-15    2
-7.86252217e+01-7.49173676e+00 8.89660986e-01 1.70119767e-02-1.13807350e-05    3
 3.88280928e-09-5.32841479e-13 1.60316121e+03 1.85001134e+01                   4
CH2OH                   C   1H   3O   1     G    300.00   3500.00 1360.00      1
 5.04534949e+00 6.02727060e-03-2.11386821e-06 3.36085906e-10-2.00987483e-14    2
-4.03584143e+03-1.57524072e+00 2.34821579e+00 1.39600168e-02-1.08632206e-05    3
 4.62498415e-09-8.08499162e-13-3.30222106e+03 1.22661977e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335655e+00 1.00905182e-02-5.12952555e-06 1.25425205e-09-1.19639106e-13    2
-1.39080170e+04 1.59916142e+01 4.32621280e+00-7.01151756e-03 3.15176939e-05    3
-3.36478617e-08 1.23454015e-11-1.43270169e+04 2.62028968e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278258e-03-2.69184211e-06 7.21357799e-10-7.43521409e-14    2
 4.05725330e+03 1.07450933e+01 4.03483979e+00-2.15836864e-03 1.18233875e-05    3
-1.18459406e-08 4.00593955e-12 3.83636392e+03 4.20008770e+00                   4
HO2CHO                  C   1H   2O   3     G    300.00   3500.00 1750.00      1
 1.00230825e+01 4.43559488e-03-1.56185338e-06 2.43413972e-10-1.38379570e-14    2
-3.81313380e+04-2.33591553e+01 2.47434345e+00 2.16898555e-02-1.63512196e-05    3
 5.87745825e-09-8.18701426e-13-3.54892793e+04 1.72835404e+01                   4
HOCHO                   H   2C   1O   2     G    200.00   3500.00 1800.00      1
 3.79473661e+00 8.42765725e-03-3.84722250e-06 8.63389842e-10-7.73674422e-14    2
-4.73118221e+04 5.12933885e+00 1.85206265e+00 1.27447105e-02-7.44476686e-06    3
 2.19581368e-09-2.62426309e-13-4.66124595e+04 1.56434956e+01                   4
OCHO                    C   1O   2H   1     G    200.00   3500.00  700.00      1
 2.58373953e+00 8.99565940e-03-4.55939788e-06 1.11902584e-09-1.07899899e-13    2
-1.67164582e+04 1.34890938e+01 4.25809175e+00-5.72067577e-04 1.59428742e-05    3
-1.84069476e-08 6.86566204e-12-1.69508675e+04 6.00851171e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959141e+00 1.57445262e-02-5.96197393e-06 1.06867182e-09-7.61012341e-14    2
-1.25948053e+04-1.43089411e+00-2.41778723e-01 2.53475709e-02-1.39645112e-05    3
 4.03257452e-09-4.87754387e-13-1.10391121e+04 2.19572625e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791360e+00 1.11042800e-02-3.71281686e-06 5.47665572e-10-2.89412605e-14    2
 1.17176215e+04-4.91382512e+00 6.75421802e-01 2.11542617e-02-1.20878017e-05    3
 3.64951180e-09-4.59753237e-13 1.33457186e+04 1.95628439e+01                   4
C2H5O2H                 C   2H   6O   2     G    300.00   3500.00 1450.00      1
 1.00876750e+01 1.40221806e-02-4.79128016e-06 7.15474136e-10-3.78163633e-14    2
-2.40669299e+04-2.56733582e+01-5.77204916e-01 4.34425389e-02-3.52261336e-05    3
 1.47085102e-08-2.45040879e-12-2.09741147e+04 2.97412031e+01                   4
C2H5O2                  C   2H   5O   2     G    300.00   3500.00 1480.00      1
 9.29919682e+00 1.29334625e-02-4.54028592e-06 7.01327864e-10-3.92078231e-14    2
-7.64002445e+03-2.14311735e+01 2.00183270e-01 3.75253910e-02-2.94645378e-05    3
 1.19284683e-08-1.93568426e-12-4.94671644e+03 2.60335034e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402718e+00 9.50595350e-03-3.15129262e-06 4.53052075e-10-2.23949160e-14    2
 3.97229102e+03-3.77420904e+00-6.02932446e-02 2.08133970e-02-1.34307867e-05    3
 4.60638300e-09-6.51687481e-13 5.51151676e+03 2.10642172e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728376e+00 7.47581589e-03-2.58984227e-06 4.05265796e-10-2.35022722e-14    2
 3.38403785e+04 1.51958752e+00 1.23421214e+00 1.56222204e-02-1.10171572e-05    3
 4.27989337e-09-6.91541508e-13 3.46967692e+04 1.68637048e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267451e+00 5.47212836e-03-2.03181547e-06 3.75019136e-10-2.77049085e-14    2
 2.58626598e+04-2.43835908e+00 7.70536982e-01 2.37107994e-02-3.66622035e-05    3
 2.95989753e-08-9.27579229e-12 2.64317975e+04 1.40907680e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788257e+00 4.21328989e-03-1.58936946e-06 2.68739191e-10-1.73346358e-14    2
 6.72874491e+04 5.32512366e+00 4.60873599e+00 1.42766785e-03 8.54158643e-07    3
-6.83903344e-10 1.21940589e-13 6.68801772e+04-1.05894068e+00                   4
C2H5OH                  C   2H   6O   1     G    300.00   3500.00 1580.00      1
 7.32490826e+00 1.39762977e-02-4.67366749e-06 6.82063686e-10-3.47025040e-14    2
-3.18909574e+04-1.38313071e+01-4.22291410e-01 3.35894614e-02-2.32937596e-05    3
 8.53864265e-09-1.27783209e-12-2.94428423e+04 2.70882146e+01                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957253e+00 2.35453826e-02-1.23415274e-05 3.08911894e-09-2.98016650e-13    2
-3.10347953e+03 1.69410914e+01 3.27852951e+00 1.44656284e-02 7.11508866e-06    3
-1.54409916e-08 6.31987996e-12-3.32593351e+03 9.84203359e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479679e+00 1.17471700e-02-4.06239752e-06 6.31554727e-10-3.61645076e-14    2
-6.24418450e+03-9.60110090e+00 1.82077786e+00 2.63431399e-02-1.89562444e-05    3
 7.38613379e-09-1.18490244e-12-4.66716293e+03 1.83437446e+01                   4
SC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1500.00      1
 6.63757422e+00 1.19924586e-02-4.07718738e-06 6.22004999e-10-3.47508086e-14    2
-9.66525354e+03-7.65007786e+00 1.23305393e+00 2.64045127e-02-1.84892415e-05    3
 7.02736238e-09-1.10231037e-12-8.04389745e+03 2.06149529e+01                   4
C2H4O2H                 C   2H   5O   2     G    300.00   3500.00 1440.00      1
 9.66417632e+00 1.29483231e-02-4.44318338e-06 6.83406485e-10-3.84804396e-14    2
 1.86599132e+03-2.38806240e+01 2.23212418e+00 3.35929124e-02-2.59479639e-05    3
 1.06393234e-08-1.76693823e-12 4.00642234e+03 1.46847780e+01                   4
C2H4O1-2                C   2H   4O   1     G    300.00   3500.00 1520.00      1
 6.04215803e+00 1.11433647e-02-3.80167463e-06 5.65226942e-10-2.94248189e-14    2
-9.44151524e+03-1.02352918e+01-2.19672856e+00 3.28246452e-02-2.51976751e-05    3
 9.94943769e-09-1.57288053e-12-6.93689371e+03 3.29622805e+01                   4
C2H3O1-2                C   2H   3O   1     G    200.00   3500.00 1800.00      1
 7.60993626e+00 6.11300596e-03-1.59366937e-06 1.28294159e-10 2.98968070e-15    2
 1.61313302e+04-1.70584528e+01 7.34197745e-02 2.28608204e-02-1.55501814e-05    3
 5.29737268e-09-7.14937891e-13 1.88444761e+04 2.37307466e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195371e+00 1.06589270e-02-3.75190329e-06 6.00731629e-10-3.66603825e-14    2
-2.30621355e+04-8.31408576e+00 9.75916637e-01 2.23167871e-02-1.34667868e-05    3
 4.19883662e-09-5.36397186e-13-2.11735621e+04 2.00785613e+01                   4
CH3CO                   C   2H   3O   1     G    300.00   3500.00 1800.00      1
 6.07689016e+00 8.12979339e-03-2.81854999e-06 4.38698308e-10-2.55171838e-14    2
-4.06801047e+03-6.15492452e+00 1.47388064e+00 1.83587034e-02-1.13426417e-05    3
 3.59576931e-09-4.63999267e-13-2.41092705e+03 1.87575232e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703792e+00 7.91358605e-03-2.83605892e-06 4.62112658e-10-2.83231300e-14    2
-1.16170812e+03-8.37157284e+00 7.37868283e-01 2.50454357e-02-2.20135026e-05    3
 1.00031294e-08-1.80836357e-12 3.76389339e+02 2.09962836e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523628e+00 6.46841658e-03-2.33588415e-06 3.83408112e-10-2.36897851e-14    2
-8.05944305e+03-4.61154401e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226118e-09-9.59140717e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420512e+00 3.89116780e-03-1.41168609e-06 2.35668534e-10-1.49424973e-14    2
 1.94026782e+04-4.94089645e+00 3.33028661e+00 1.20351629e-02-1.14247949e-05    3
 5.70731267e-09-1.13618105e-12 2.00087543e+04 7.53650387e+00                   4
HCOOH                   C   1H   2O   2     G    300.00   3500.00 1640.00      1
 5.21581644e+00 5.48253641e-03-1.72756112e-06 2.25438491e-10-8.81949923e-15    2
-4.56198641e+04-2.59494559e+00 1.19691275e+00 1.52847405e-02-1.06929917e-05    3
 3.86992247e-09-5.64381081e-13-4.43016637e+04 1.87820781e+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   3500.00 1760.00      1
 1.40469381e+01 2.48483420e-03 1.65900438e-06-8.55133987e-10 9.82287243e-14    2
-2.73756816e+04-4.36816972e+01 2.64892548e+00 2.83894083e-02-2.04187576e-05    3
 7.50765465e-09-1.08966739e-12-2.33635811e+04 1.77505788e+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772146e-02-4.04888400e-06 6.94756703e-10-4.56573678e-14    2
-7.51809422e+04-3.74730275e+01-2.33886891e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164714e-12-7.15304886e+04 3.67067395e+01                   4
CH3OCHO                 C   2H   4O   2     G    300.00   3500.00  700.00      1
 5.02910661e+00-2.87377520e-02 6.15808971e-05-2.98073518e-08 4.29774802e-12    2
-4.07046731e+04 1.82412179e+01 4.01576605e-08-2.13669220e-10 3.62011546e-13    3
 2.88411213e-08-1.66481352e-11-4.00005982e+04 4.07099937e+01                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849389e-09-3.11411020e-13    2
-2.07588781e+04 1.60124236e+01 4.66126892e+00 9.68655559e-03 1.14715527e-05    3
-1.83003964e-08 7.03409935e-12-2.10634335e+04 6.60518521e+00                   4
CH2OHCHO                C   2H   4O   2     G    300.00   3500.00 1800.00      1
 8.91045186e+00 9.14305837e-03-2.53718677e-06 2.39203913e-10 8.50819808e-16    2
-4.09945450e+04-1.84179622e+01 1.56305396e+00 2.54706093e-02-1.61434792e-05    3
 5.27857147e-09-6.99061341e-13-3.83494818e+04 2.13476880e+01                   4
CHOCHO                  C   2H   2O   2     G    300.00   3500.00 1570.00      1
 9.97760258e+00 4.26981224e-03-1.12729433e-06 7.37809077e-11 5.98360554e-15    2
-2.96900177e+04-2.75230973e+01 7.08345766e-01 2.78857532e-02-2.36902952e-05    3
 9.65467301e-09-1.51963616e-12-2.67794711e+04 2.13768445e+01                   4
O2C2H4O2H               C   2H   5O   4     G    300.00   3500.00 1800.00      1
 1.24323243e+01 1.62358927e-02-6.84260319e-06 1.39267431e-09-1.12911127e-13    2
-1.87641105e+04-2.90906767e+01 5.81911522e+00 3.09319128e-02-1.90892866e-05    3
 5.92848300e-09-7.42884555e-13-1.63833552e+04 6.70139036e+00                   4
HO2CH2CHO               C   2H   4O   3     G    300.00   3500.00 1240.00      1
 1.23807018e+01 1.08772146e-02-4.04888400e-06 6.94756703e-10-4.56573678e-14    2
-7.51809422e+04-3.74730275e+01-2.33886891e+00 5.83597007e-02-6.14873753e-05    3
 3.15756660e-08-6.27164714e-12-7.15304886e+04 3.67067395e+01                   4
C3H8                    C   3H   8          G    300.00   3500.00 1690.00      1
 8.33847007e+00 1.79340922e-02-5.80534982e-06 7.91037710e-10-3.43401229e-14    2
-1.70816233e+04-2.27461799e+01-1.38651265e+00 4.09518028e-02-2.62352705e-05    3
 8.85017800e-09-1.22652064e-12-1.37945792e+04 2.92742161e+01                   4
IC3H7                   C   3H   7          G    300.00   3500.00 1800.00      1
 6.05951250e+00 1.82035621e-02-6.54041321e-06 1.09272144e-09-7.13189355e-14    2
 7.29671818e+03-6.80793081e+00-6.08211221e-01 3.30207259e-02-1.88880497e-05    3
 5.66592015e-09-7.06485423e-13 9.69709872e+03 2.92791809e+01                   4
NC3H7                   C   3H   7          G    300.00   3500.00 1590.00      1
 7.21724981e+00 1.65877265e-02-5.58902439e-06 8.31338517e-10-4.40999327e-14    2
 8.50975634e+03-1.26938766e+01-1.37086177e-01 3.50892007e-02-2.30432453e-05    3
 8.14967014e-09-1.19478101e-12 1.08484352e+04 2.61969991e+01                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755201e+00 1.65820017e-02-6.59972302e-06 1.29512916e-09-1.03784375e-13    2
-3.79456071e+02-1.05616188e+01-8.55987190e-02 3.08112255e-02-1.84574096e-05    3
 5.68686491e-09-7.13747674e-13 1.92567819e+03 2.40935688e+01                   4
C3H5-A                  C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877792e+00 1.04611885e-02-3.15379708e-06 3.85306883e-10-1.26413688e-14    2
 1.71766363e+04-2.28181758e+01-3.57888096e-01 3.27028536e-02-2.40053581e-05    3
 9.07345729e-09-1.37016487e-12 2.00235695e+04 2.42845603e+01                   4
C3H5-S                  C   3H   5          G    300.00   3500.00 1800.00      1
 6.52599516e+00 1.37686655e-02-5.50691342e-06 1.07278366e-09-8.39560018e-14    2
 2.86430050e+04-9.99635699e+00 1.54227621e+00 2.48435965e-02-1.47360226e-05    3
 4.49097224e-09-5.58704416e-13 3.04371438e+04 1.69765696e+01                   4
C3H5-T                  C   3H   5          G    300.00   3500.00  770.00      1
 1.49331935e+00 2.33788729e-02-1.18550710e-05 2.86552469e-09-2.68203790e-13    2
 2.87117775e+04 1.76892214e+01 2.52238868e+00 1.80330582e-02-1.44114628e-06    3
-6.15086038e-09 2.65919396e-12 2.85533009e+04 1.29935192e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079978e+00 1.37589660e-02-5.15319199e-06 9.32421983e-10-6.74695911e-14    2
 7.77376170e+03-2.10036658e+01 9.27196847e-01 3.40908988e-02-2.40959865e-05    3
 8.77622923e-09-1.28545208e-12 1.04088818e+04 2.23747992e+01                   4
C3H6O                   C   3H   6O   1     G    300.00   3500.00 1550.00      1
 9.00938221e+00 1.57632590e-02-5.29374356e-06 7.64253420e-10-3.74126441e-14    2
-1.56669515e+04-2.44960178e+01-1.88321637e+00 4.38731909e-02-3.24969034e-05    3
 1.24645372e-08-1.92455519e-12-1.22902459e+04 3.28282089e+01                   4
CH3CHCHO                C   3H   5O   1     G    300.00   3500.00 1800.00      1
 6.70347362e+00 1.89922318e-02-9.18109976e-06 2.14445657e-09-1.96154637e-13    2
-6.21094363e+03-1.05801331e+01 2.92067498e-01 3.32398010e-02-2.10540741e-05    3
 6.54185446e-09-8.06904344e-13-3.90283743e+03 2.41197343e+01                   4
AC4H7OOH                C   4H   8O   2     G    300.00   3500.00 1660.00      1
 1.22738272e+01 2.55483383e-02-9.81265076e-06 1.82078670e-09-1.35039880e-13    2
-1.24525960e+04-3.36837474e+01 1.60151447e+00 5.12647544e-02-3.30503762e-05    3
 1.11532065e-08-1.54052480e-12-8.90938817e+03 2.32129081e+01                   4
CH3CHCO                 C   3H   4O   1     G    300.00   3500.00 1280.00      1
 6.99681463e+00 1.49445085e-02-6.71568578e-06 1.45955079e-09-1.25293200e-13    2
-1.29366480e+04-1.07908059e+01 1.50068776e+00 3.21199049e-02-2.68431035e-05    3
 1.19425809e-08-2.17276001e-12-1.15296395e+04 1.70816035e+01                   4
AC3H5OOH                C   3H   6O   2     G    298.00   3500.00 1800.00      1
 1.36957657e+01 1.27112963e-02-4.21186263e-06 6.49030109e-10-3.94931201e-14    2
-1.11479407e+04-4.31791017e+01 4.22354618e+00 3.37606729e-02-2.17530098e-05    3
 7.14575129e-09-9.41815506e-13-7.73794171e+03 8.08652617e+00                   4
C3H6OH1-2               C   3H   7O   1     G    300.00   3500.00 1800.00      1
 8.46016352e+00 1.89669003e-02-7.38013554e-06 1.39189577e-09-1.05413394e-13    2
-1.21581707e+04-1.51603325e+01 4.08605477e-01 3.68592515e-02-2.22904282e-05    3
 6.91422639e-09-8.72403758e-13-9.25960980e+03 2.84163793e+01                   4
C3H6OH2-1               C   3H   7O   1     G    300.00   3500.00 1590.00      1
 8.99548234e+00 1.75103792e-02-6.94615357e-06 1.37004323e-09-1.07539337e-13    2
-1.65436320e+04-1.93287236e+01 1.31207693e+00 3.68397010e-02-2.51813628e-05    3
 9.01583327e-09-1.30970758e-12-1.41003090e+04 2.13023225e+01                   4
HOC3H6O2                C   3H   7O   3     G    300.00   3500.00 1480.00      1
 1.24409055e+01 2.15172909e-02-8.97737594e-06 1.82414691e-09-1.48047122e-13    2
-3.10315628e+04-3.23089026e+01 2.93449048e+00 4.72103044e-02-3.50175923e-05    3
 1.35539741e-08-2.12943685e-12-2.82176640e+04 1.72809693e+01                   4
SC3H5OH                 C   3H   6O   1     G    300.00   3500.00 1260.00      1
 7.83167544e+00 1.85990426e-02-7.98421837e-06 1.67672191e-09-1.40411942e-13    2
-2.22362405e+04-1.56369776e+01-5.71229655e-02 4.36428470e-02-3.77982713e-05    3
 1.74513531e-08-3.27029908e-12-2.02482633e+04 2.42451083e+01                   4
C3H5OH                  C   3H   6O   1     G    300.00   3500.00 1630.00      1
 9.39463114e+00 1.51343106e-02-4.86246277e-06 6.64177251e-10-2.94552533e-14    2
-2.20582199e+04-2.45922026e+01 4.73537668e-01 3.70265645e-02-2.50087087e-05    3
 8.90395064e-09-1.29322418e-12-1.91499434e+04 2.28055845e+01                   4
CH2CCH2OH               C   3H   5O   1     G    300.00   3500.00 1800.00      1
 7.15397365e+00 1.62590933e-02-7.06959971e-06 1.52062107e-09-1.30983749e-13    2
 1.01359982e+04-8.36739478e+00 2.39300609e+00 2.68390212e-02-1.58862063e-05    3
 4.78603091e-09-5.84512894e-13 1.18499465e+04 1.73999548e+01                   4
C3H4-P                  C   3H   4          G    300.00   3500.00 1570.00      1
 6.45797858e+00 1.06371316e-02-3.61161722e-06 5.39412692e-10-2.85851276e-14    2
 1.94136786e+04-1.10770989e+01 1.72714322e+00 2.26902153e-02-1.51273023e-05    3
 5.42930020e-09-8.07229635e-13 2.08991609e+04 1.38804115e+01                   4
C3H4-A                  C   3H   4          G    300.00   3500.00 1420.00      1
 6.37608366e+00 1.10282079e-02-3.89476312e-06 6.16686075e-10-3.59564767e-14    2
 2.00917847e+04-1.13283006e+01 5.08248695e-01 2.75573205e-02-2.13550933e-05    3
 8.81402419e-09-1.47914981e-12 2.17582498e+04 1.90382079e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057760e+00 1.05635748e-02-4.84060957e-06 1.09040070e-09-9.80036150e-14    2
 4.00565408e+04-5.04125047e+00 1.75584152e+00 2.95861275e-02-3.88094537e-05    3
 2.80498008e-08-8.12163460e-12 4.07276565e+04 1.35345461e+01                   4
C3H2                    C   3H   2          G    300.00   3500.00 1260.00      1
 6.42043188e+00 6.05128867e-03-2.30888142e-06 4.10631877e-10-2.84293477e-14    2
 6.08598164e+04-8.32404332e+00 2.15397882e+00 1.95955841e-02-1.84330427e-05    3
 8.94193412e-09-1.72114805e-12 6.19349626e+04 1.32451538e+01                   4
C3H3O                   H   3C   3O   1     G    298.15   3500.00  860.00      1
 4.35781247e+00 1.92087074e-02-1.19701078e-05 3.82443985e-09-4.99532170e-13    2
 3.14370432e+04 4.14502711e+00 7.87593033e-01 3.58143792e-02-4.09334889e-05    3
 2.62766733e-08-7.02634421e-12 3.20511210e+04 2.08308013e+01                   4
C2H5CHO                 C   3H   6O   1     G    300.00   3500.00 1710.00      1
 9.33264603e+00 1.46861072e-02-4.56011956e-06 5.69518137e-10-1.90908111e-14    2
-2.69164882e+04-2.52385565e+01-9.86882745e-02 3.67477079e-02-2.39124009e-05    3
 8.11426720e-09-1.12212430e-12-2.36909719e+04 2.53220280e+01                   4
CH2CH2CHO               C   3H   5O   1     G    300.00   3500.00  700.00      1
 1.38640400e+00 2.84363938e-02-1.56688640e-05 4.07196321e-09-4.03232083e-13    2
 6.14151634e+02 2.19844218e+01 2.41071832e+00 2.25831692e-02-3.12623980e-06    3
-7.87339320e-09 3.86296664e-12 4.70747631e+02 1.74080446e+01                   4
RALD3BG                 C   3H   5O   1     G    300.00   3500.00 1140.00      1
-6.08013768e+00 4.60180077e-02-2.61696720e-05 6.65382129e-09-6.35305356e-13    2
-2.14966002e+03 5.90959839e+01 7.04072885e+00-2.01204289e-05 3.44068124e-05    3
-2.87710234e-08 7.13330094e-12-5.14121758e+03-5.92381683e+00                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597838e+00 1.12038372e-02-3.67974366e-06 5.08180254e-10-2.25803378e-14    2
-1.23719484e+04-2.08137560e+01 8.18908044e-01 3.22215131e-02-2.33838148e-05    3
 8.71820988e-09-1.30539747e-12-9.68168587e+03 2.36968522e+01                   4
CH3COCH3                C   3H   6O   1     G    300.00   3500.00 1790.00      1
 9.79507855e+00 1.35932466e-02-4.01642284e-06 4.43034307e-10-7.94380264e-15    2
-3.07542949e+04-2.70699391e+01-7.54581319e-03 3.54985524e-02-2.23728244e-05    3
 7.27968292e-09-9.62782995e-13-2.72449554e+04 2.59292980e+01                   4
CH3COCH2                C   3H   5O   1     G    300.00   3500.00 1590.00      1
 8.40473847e+00 1.29432044e-02-4.25667367e-06 6.02254913e-10-2.86748420e-14    2
-7.89528923e+03-1.63899805e+01 1.00367440e+00 3.15622335e-02-2.18217955e-05    3
 7.96708585e-09-1.18666713e-12-5.54175085e+03 2.27480006e+01                   4
NC4H10                  C   4H  10          G    300.00   3500.00 1800.00      1
 1.54355362e+01 1.56272553e-02-3.14852000e-06-5.94424183e-11 5.32964635e-14    2
-2.28455262e+04-6.02417835e+01-1.20836758e+00 5.26137081e-02-3.39705640e-05    3
 1.13561294e-08-1.53219963e-12-1.68537208e+04 2.98384958e+01                   4
PC4H9                   C   4H   9          G    300.00   3500.00  950.00      1
 3.94763005e+00 3.16286394e-02-1.12984867e-05 1.11637451e-09 5.54031595e-14    2
 6.05554723e+03 7.76350068e+00-2.76188368e-01 4.94131380e-02-3.93792740e-05    3
 2.08221901e-08-5.13033779e-12 6.85807273e+03 2.79243294e+01                   4
SC4H9                   C   4H   9          G    300.00   3500.00  850.00      1
 3.40122925e+00 3.20901864e-02-1.12255471e-05 9.71712126e-10 8.30726255e-14    2
 4.66283102e+03 1.05291640e+01 2.36336467e-01 4.69837995e-02-3.75083938e-05    3
 2.15857095e-08-5.97986778e-12 5.20086279e+03 2.52835872e+01                   4
IC4H10                  C   4H  10          G    300.00   3500.00 1260.00      1
 5.51955794e+00 3.23747266e-02-1.18655436e-05 1.37455178e-09 1.57073476e-14    2
-1.97025810e+04-6.34483422e+00-1.85965328e+00 5.58007940e-02-3.97537190e-05    3
 1.61302002e-08-2.91200067e-12-1.78430198e+04 3.09610166e+01                   4
IC4H9                   C   4H   9          G    300.00   3500.00 1430.00      1
 7.95880517e+00 2.55088283e-02-8.62221491e-06 8.09648923e-10 4.02033219e-14    2
 3.37759298e+03-1.61084037e+01-1.15582376e+00 5.10042938e-02-3.53657102e-05    3
 1.32774789e-08-2.13948724e-12 5.98437685e+03 3.11244820e+01                   4
TC4H9                   C   4H   9          G    300.00   3500.00 1400.00      1
 7.90871688e+00 2.55264450e-02-8.65284050e-06 8.24419703e-10 3.80550654e-14    2
 8.35470581e+02-1.73299272e+01-1.29900233e+00 5.18342142e-02-3.68397360e-05    3
 1.42467509e-08-2.35878979e-12 3.41363196e+03 3.01901373e+01                   4
IC4H8                   C   4H   8          G    300.00   3500.00 1800.00      1
 7.63433967e+00 2.47722696e-02-1.05415828e-05 2.18152373e-09-1.80119594e-13    2
-6.21385767e+03-1.72949366e+01 7.17301598e-01 4.01434653e-02-2.33509125e-05    3
 6.92571993e-09-8.39035733e-13-3.72372397e+03 2.01415164e+01                   4
IC4H7                   C   4H   7          G    300.00   3500.00  700.00      1
 1.18177119e+00 3.67769036e-02-1.77031336e-05 3.74786264e-09-2.92191282e-13    2
 1.31214242e+04 2.00120539e+01 3.86129999e+00 2.14653105e-02 1.51074231e-05    3
-2.75002866e-08 1.08678620e-11 1.27462902e+04 8.04059711e+00                   4
IC4H7O                  C   4H   7O   1     G    300.00   3500.00 1800.00      1
 1.18822163e+01 1.89918532e-02-7.42296498e-06 1.41442848e-09-1.08683660e-13    2
 1.15971319e+03-3.56333819e+01 1.50010972e+00 4.20632012e-02-2.66490883e-05    3
 8.53521488e-09-1.09768177e-12 4.89727156e+03 2.05567447e+01                   4
C4H8-1                  C   4H   8          G    300.00   3500.00 1800.00      1
 1.03330449e+01 1.99470428e-02-7.40538998e-06 1.30472507e-09-9.09598189e-14    2
-5.56551437e+03-3.07722296e+01-6.91489887e-01 4.44460090e-02-2.78211951e-05    3
 8.86613439e-09-1.14115556e-12-1.59668184e+03 2.88948525e+01                   4
C4H8-2                  C   4H   8          G    300.00   3500.00 1800.00      1
 5.15907399e+00 2.89997694e-02-1.32974598e-05 2.96139017e-09-2.60424474e-13    2
-4.76704683e+03-3.39008062e+00 5.60608454e-01 3.92185817e-02-2.18131368e-05    3
 6.11534459e-09-6.98473698e-13-3.11159924e+03 2.14977742e+01                   4
C4H71-3                 C   4H   7          G    300.00   3500.00 1420.00      1
 8.33017753e+00 1.98466503e-02-6.37614062e-06 5.28652771e-10 3.81103731e-14    2
 1.19533850e+04-1.83767118e+01-1.12550124e+00 4.64823652e-02-3.45124591e-05    3
 1.37381920e-08-2.28751273e-12 1.46387978e+04 3.05571711e+01                   4
C4H71-4                 C   4H   7          G    300.00   3500.00 1530.00      1
 8.45916998e+00 1.93968541e-02-5.99075606e-06 3.82147973e-10 5.73994806e-14    2
 1.98988324e+04-1.80212793e+01-3.29329051e-01 4.23733221e-02-2.85167051e-05    3
 1.01973763e-08-1.54639600e-12 2.25881131e+04 2.81156134e+01                   4
C4H71-O                 C   4H   7O   1     G    300.00   3500.00 1600.00      1
 1.37371777e+01 1.70982846e-02-6.55972543e-06 1.21466090e-09-8.98269615e-14    2
-3.28789073e+01-4.64105970e+01-1.48200925e+00 5.51462520e-02-4.22296948e-05    3
 1.60771481e-08-2.41209059e-12 4.83726091e+03 3.41662556e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872521e+00 1.50139591e-02-5.06688177e-06 7.84148096e-10-4.70262839e-14    2
 8.60829987e+03-2.47389586e+01 4.65225109e-01 3.46661815e-02-2.14437338e-05    3
 6.84964885e-09-8.89456944e-13 1.17919599e+04 2.31239087e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794385e-03 4.88814513e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742307e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777119e+00 1.26498258e-02-4.62248952e-06 7.81217086e-10-5.07629111e-14    2
 3.13366016e+04-1.49692661e+01 7.13119719e-01 3.41836288e-02-2.96617953e-05    3
 1.37214268e-08-2.55855549e-12 3.31283217e+04 2.03030643e+01                   4
C4H3                    C   4H   3          G    300.00   3500.00 1590.00      1
 1.30208969e+01 1.53590365e-03 1.80568199e-06-9.30237202e-10 1.18077197e-13    2
 6.01811751e+04-4.25791500e+01 2.34662667e+00 2.83894138e-02-2.35278181e-05    3
 9.69177542e-09-1.55205057e-12 6.35755930e+04 1.38680560e+01                   4
C4H2                    C   4H   2          G    300.00   3500.00  720.00      1
 7.13414724e+00 1.00526311e-02-4.84819229e-06 1.14884612e-09-1.07722844e-13    2
 5.27577825e+04-1.36443510e+01-4.34753652e-01 5.21020805e-02-9.24512119e-05    3
 8.22627532e-08-2.82722739e-11 5.38477042e+04 2.03848058e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055544e+01 1.99961046e-02-7.07935462e-06 1.10673029e-09-6.24178906e-14    2
 4.11452291e+03-4.24445090e+01-6.99882110e+00 7.24907868e-02-6.29247613e-05    3
 2.75111779e-08-4.74405754e-12 9.33275680e+03 5.31863191e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152220e+01 1.47750067e-02-3.90939181e-06 2.82308156e-10 1.62511622e-14    2
 1.91167581e+04-5.54965184e+01-3.67012639e+00 6.11476948e-02-4.84985149e-05    3
 1.93374890e-08-3.03746371e-12 2.47593868e+04 3.97971310e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331261e+01 1.77269650e-02-6.33615685e-06 1.00236866e-09-5.75481757e-14    2
 3.49856300e+04-3.80075864e+01-6.76261385e+00 6.95132669e-02-6.22206553e-05    3
 2.78054854e-08-4.87825263e-12 3.99884457e+04 5.47375207e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786764e+01 1.28174257e-02-3.11961936e-06 1.29368392e-10 2.76958521e-14    2
 9.43770579e+03-5.26289052e+01-4.05866643e+00 5.60992486e-02-4.29495178e-05    3
 1.64197154e-08-2.47082363e-12 1.51874796e+04 4.10783319e+01                   4
C5H5                    C   5H   5          G    300.00   3500.00  700.00      1
 4.01652580e+00 2.68451889e-02-1.26423017e-05 2.78092329e-09-2.35299432e-13    2
 2.91110159e+04 1.44025771e+00-2.58737429e+00 6.45817609e-02-9.35063844e-05    3
 7.97943354e-08-2.77400895e-11 3.00355619e+04 3.09448125e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1800.00      1
-1.21144532e+02 2.92206047e-01-1.95445890e-04 5.59670212e-08-5.79656630e-12    2
 5.40571659e+04 6.85330239e+02 7.45334840e+00 6.43297952e-03 4.26983328e-05    3
-3.22345427e-08 6.45365091e-12 7.76192901e+03-1.06683155e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248658e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987877e+01                   4
NC5H12                  C   5H  12          G    300.00   3500.00 1800.00      1
 2.12559082e+01 1.49866375e-02-1.56738312e-06-4.84518435e-10 9.00436509e-14    2
-2.80668702e+04-9.05497671e+01-1.97000865e+00 6.65997861e-02-4.45783403e-05    3
 1.54454657e-08-2.12245414e-12-1.97055401e+04 3.51537401e+01                   4
NC5H11                  C   5H  11          G    300.00   3500.00 1800.00      1
 6.93193785e+00 3.75440987e-02-1.65478566e-05 3.53633643e-09-2.99976701e-13    2
-1.73087074e+03-8.88710672e+00-3.57520449e+00 6.08933039e-02-3.60055276e-05    3
 1.07428812e-08-1.30088570e-12 2.05170050e+03 4.79797395e+01                   4
NEOC5H12                C   5H  12          G    300.00   3500.00 1700.00      1
 1.58220811e+01 2.73824077e-02-1.01392581e-05 1.77707009e-09-1.22756971e-13    2
-2.85197010e+04-6.62488521e+01-2.62463460e+00 7.07864446e-02-4.84369376e-05    3
 1.67957680e-08-2.33138901e-12-2.22478177e+04 3.25342362e+01                   4
NEOC5H11                C   5H  11          G    300.00   3500.00 1670.00      1
 1.43276289e+01 2.66845577e-02-1.02158264e-05 1.86929104e-09-1.35803312e-13    2
-2.94216421e+03-5.15145769e+01-1.29689709e+00 6.41085720e-02-4.38302105e-05    3
 1.52882069e-08-2.14462305e-12 2.27642747e+03 3.18773552e+01                   4
NC5H10                  C   5H  10          G    300.00   3500.00 1800.00      1
 1.11929736e+01 2.82582223e-02-1.13863841e-05 2.22526491e-09-1.74280993e-13    2
-1.02483443e+04-3.39253533e+01-6.89551964e-01 5.46638348e-02-3.33910611e-05    3
 1.03751453e-08-1.30620882e-12-5.97063504e+03 3.03853541e+01                   4
NC5H9-3                 C   5H   9          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
B1M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.21299340e+01 2.65376145e-02-1.02995525e-05 1.93064538e-09-1.45051208e-13    2
-1.11266091e+04-3.96207198e+01-6.39002025e-01 5.49130280e-02-3.39457304e-05    3
 1.06884890e-08-1.36141838e-12-6.52979211e+03 2.94874259e+01                   4
B1M3                    C   5H  10          G    300.00   3500.00 1800.00      1
 1.31681365e+01 2.49963287e-02-9.30063098e-06 1.64277853e-09-1.14892348e-13    2
-1.09953810e+04-4.60629132e+01-8.44094903e-01 5.61346208e-02-3.52492077e-05    3
 1.12533625e-08-1.44969568e-12-5.95097767e+03 2.97742066e+01                   4
B2M2                    C   5H  10          G    300.00   3500.00 1800.00      1
 9.73411699e+00 3.08235227e-02-1.30972997e-05 2.71635425e-09-2.25270435e-13    2
-1.14704814e+04-2.74877025e+01 1.14407401e-01 5.22006552e-02-3.09115767e-05    3
 9.31423462e-09-1.14164271e-12-8.00738598e+03 2.45761726e+01                   4
CYC5H8                  C   5H   8          G    300.00   3500.00 1460.00      1
 8.43099915e+00 2.71082714e-02-1.07932862e-05 1.95387666e-09-1.31111174e-13    2
-1.09862538e+03-2.37608447e+01-6.56863980e+00 6.82031726e-02-5.30140751e-05    3
 2.12327757e-08-3.43229252e-12 3.28126920e+03 5.42801525e+01                   4
C5H7                    C   5H   7          G    300.00   3500.00 1430.00      1
 7.72404525e+00 2.56072196e-02-8.76350316e-06 8.66193959e-10 3.30416650e-14    2
 2.30808142e+04-1.69352935e+01 2.31765047e-01 4.65646468e-02-3.07468184e-05    3
 1.11148258e-08-1.75867718e-12 2.52236063e+04 2.18904247e+01                   4
LC5H8                   C   5H   8          G    300.00   3500.00 1430.00      1
 8.95829159e+00 2.51033002e-02-8.43679234e-06 8.19905621e-10 3.11426511e-14    2
 4.67953300e+03-2.40439628e+01 1.19183502e+00 4.68276543e-02-3.12245763e-05    3
 1.14435811e-08-1.82614328e-12 6.90073958e+03 1.62025638e+01                   4
DIALLYL                 C   6H  10          G    300.00   3500.00 1670.00      1
 1.46885479e+01 2.58341295e-02-9.34005191e-06 1.60362033e-09-1.08722036e-13    2
 2.72208305e+03-5.11904320e+01-8.93391061e-01 6.31561390e-02-4.28628149e-05    3
 1.49859609e-08-2.11206643e-12 7.92645066e+03 3.19742027e+01                   4
RC6H9A                  C   6H   9          G    300.00   3500.00 1310.00      1
 1.02179198e+01 3.31131696e-02-1.50182299e-05 3.28859653e-09-2.83959224e-13    2
 2.30740211e+04-2.53806643e+01-2.61882183e+00 7.23093274e-02-5.98993266e-05    3
 2.61288493e-08-4.64278609e-12 2.64372474e+04 4.00154625e+01                   4
CYC6H8                  C   6H   8          G    300.00   3500.00 1490.00      1
 8.66772261e+00 3.45074855e-02-1.63846780e-05 3.69260974e-09-3.24421025e-13    2
 5.74022138e+03-2.73566208e+01-6.91358136e+00 7.63364895e-02-5.84944135e-05    3
 2.25336547e-08-3.48567018e-12 1.03834500e+04 5.40276160e+01                   4
CYC6H10                 C   6H  10          G    300.00   3500.00 1800.00      1
 1.51624858e+01 2.76360017e-02-1.05259858e-05 1.89586361e-09-1.35054773e-13    2
-9.29985245e+03-6.25064559e+01-6.01517655e+00 7.46974737e-02-4.97438791e-05    3
 1.64210093e-08-2.15243611e-12-1.67589399e+03 5.21114707e+01                   4
RCYC6H9                 C   6H   9          G    300.00   3500.00 1800.00      1
 1.41670463e+01 2.75651338e-02-1.13337615e-05 2.23021652e-09-1.74683445e-13    2
 7.93866332e+03-5.85441979e+01-6.48639356e+00 7.34616669e-02-4.95808724e-05    3
 1.63958131e-08-2.14212742e-12 1.53739017e+04 5.32365273e+01                   4
CYC6H12                 C   6H  12          G    300.00   3500.00 1800.00      1
 1.12578097e+01 4.34354098e-02-2.02455774e-05 4.54245292e-09-4.01195170e-13    2
-2.30439963e+04-4.47863376e+01-9.43363126e+00 8.94163897e-02-5.85630607e-05    3
 1.87341134e-08-2.37225913e-12-1.55950776e+04 6.72000574e+01                   4
CYC6H11                 C   6H  11          G    300.00   3500.00 1800.00      1
 1.12879190e+01 3.94798364e-02-1.80474738e-05 3.97976999e-09-3.47933573e-13    2
 4.69934406e+02-4.15743644e+01-9.20200373e+00 8.50129981e-02-5.59917752e-05    3
 1.80332150e-08-2.29980093e-12 7.84630661e+03 6.93213721e+01                   4
NC6H12                  C   6H  12          G    300.00   3500.00 1780.00      1
 2.80951654e+01 5.24635942e-03 6.43208138e-06-3.19131389e-09 4.01093698e-13    2
-1.79767847e+04-1.24497292e+02-1.85358315e+00 7.25469181e-02-5.02818725e-05    3
 1.80498673e-08-2.58221827e-12-7.31503024e+03 3.72569567e+01                   4
NC7H16                  C   7H  16          G    300.00   3500.00 1800.00      1
 3.10696120e+01 1.73458864e-02-4.57663884e-07-1.06280964e-09 1.59098857e-13    2
-3.76541592e+04-1.40920497e+02-2.76912812e+00 9.25430866e-02-6.31219974e-05    3
 2.21462028e-08-3.06437509e-12-2.54722127e+04 4.22218230e+01                   4
NC7H15                  C   7H  15          G    300.00   3500.00 1800.00      1
 1.58938298e+01 4.32851195e-02-1.83429598e-05 3.81524632e-09-3.18291961e-13    2
-8.33589206e+03-5.34387877e+01-1.03213606e+00 8.08983770e-02-4.96873411e-05    3
 1.54242764e-08-1.93065725e-12-2.24254435e+03 3.81680705e+01                   4
NC7H14                  C   7H  14          G    300.00   3500.00 1800.00      1
 1.82668105e+01 3.59607889e-02-1.37346402e-05 2.52229049e-09-1.85248240e-13    2
-1.87497345e+04-6.92309266e+01-1.22797309e+00 7.92825302e-02-4.98360912e-05    3
 1.58931983e-08-2.04231877e-12-1.17316124e+04 3.62789089e+01                   4
NC7H13                  C   7H  13          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
IC8H18                  C   8H  18          G    300.00   3500.00 1390.00      1
 2.06155885e+01 4.43694094e-02-1.35968858e-05 1.75327622e-09-6.83090879e-14    2
-3.76580614e+04-8.42148793e+01-5.96912081e+00 1.20872170e-01-9.61538217e-05    3
 4.13489289e-08-7.18982936e-12-3.02675122e+04 5.27954202e+01                   4
IC8H17                  C   8H  17          G    300.00   3500.00 1530.00      1
 2.65104230e+01 3.01796816e-02-5.82184990e-06 1.42085851e-11 7.60110760e-14    2
-1.80373025e+04-1.14981197e+02-3.32961207e+00 1.08192845e-01-8.23053435e-05    3
 3.33403496e-08-5.36943680e-12-8.90625182e+03 4.16697269e+01                   4
IC8H16                  C   8H  16          G    300.00   3500.00 1400.00      1
 1.88616063e+01 4.14292819e-02-1.28170544e-05 1.66806735e-09-6.58961709e-14    2
-2.24684067e+04-7.38514296e+01-5.35586581e+00 1.10622059e-01-8.69521729e-05    3
 3.69705048e-08-6.36990285e-12-1.56875145e+04 5.11323811e+01                   4
DIMEPTD                 C   7H  12          G    300.00   3500.00 1310.00      1
 1.53755546e+01 3.27318283e-02-1.05955708e-05 1.52102630e-09-7.69415912e-14    2
-6.19682930e+03-5.37226046e+01-1.29247813e+00 8.36265847e-02-6.88720094e-05    3
 3.11782470e-08-5.73671653e-12-1.82980473e+03 3.11918393e+01                   4
C7H8                    C   7H   8          G    200.00   3500.00 1740.00      1
 1.92535108e+01 1.64137602e-02-3.61135948e-06 2.27424888e-11 5.04456794e-14    2
-3.67626229e+03-8.27561068e+01-4.42382865e+00 7.08444256e-02-5.05343469e-05    3
 1.80008986e-08-2.53262272e-12 4.56345183e+03 4.45878951e+01                   4
C7H7                    C   7H   7          G    200.00   3500.00 1600.00      1
 1.77148781e+01 1.72901839e-02-4.74309316e-06 3.88421745e-10 1.27959347e-14    2
 1.68881058e+04-7.24712964e+01-3.23806381e+00 6.96725387e-02-5.38515508e-05    3
 2.08502791e-08-3.18436927e-12 2.35930472e+04 3.84624951e+01                   4
CH3C6H4                 C   7H   7          G    200.00   3500.00 1730.00      1
 1.83842182e+01 1.52647348e-02-3.43004338e-06 5.73661648e-11 4.21798063e-14    2
 2.84624024e+04-7.44700925e+01-2.82564598e+00 6.43048832e-02-4.59504033e-05    3
 1.64428613e-08-2.32566631e-12 3.58010154e+04 3.94808224e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1330.00      1
 1.39867712e+01 2.02277643e-02-7.36599500e-06 1.21196288e-09-7.46105017e-14    2
-1.80542263e+04-5.08485811e+01-5.47325435e+00 7.87541571e-02-7.33732049e-05    3
 3.42982836e-08-6.29384373e-12-1.28778595e+04 4.85843830e+01                   4
C6H5O                   C   6H   5O   1     G    300.00   3500.00 1320.00      1
 1.34428169e+01 1.79658729e-02-6.67332779e-06 1.12237517e-09-7.10809501e-14    2
 4.07683819e+02-4.72500520e+01-4.80707078e+00 7.32685627e-02-6.95172935e-05    3
 3.28617518e-08-6.08232652e-12 5.22565416e+03 4.58618544e+01                   4
C6H5CHO                 C   7H   6O   1     G    200.00   3500.00 1630.00      1
 2.06104936e+01 1.34209230e-02-2.83635978e-06-5.48103783e-11 5.23167108e-14    2
-1.43315560e+04-8.70895599e+01-3.50845143e+00 7.26085180e-02-5.73034718e-05    3
 2.22221271e-08-3.36439149e-12-6.46877992e+03 4.10544422e+01                   4
C7H6                    C   7H   6          G    300.00   3500.00 1290.00      1
 1.11282362e+01 2.73165807e-02-1.25329645e-05 2.76951413e-09-2.40721375e-13    2
 3.69620905e+04-3.50553513e+01-3.97785296e+00 7.41571673e-02-6.69987629e-05    3
 3.09172135e-08-5.69570188e-12 4.08594615e+04 4.16694449e+01                   4
C7H5                    C   7H   5          G    300.00   3500.00 1250.00      1
 1.21079560e+01 2.22665290e-02-9.87308080e-06 2.11666746e-09-1.79360812e-13    2
 5.15977924e+04-3.78517160e+01-2.81419579e+00 7.00174146e-02-6.71741435e-05    3
 3.26772342e-08-6.29147417e-12 5.53283304e+04 3.74688223e+01                   4
CYC5H4                  C   5H   4          G    200.00   3500.00 1310.00      1
 6.52292919e+00 1.75112106e-02-7.24525264e-06 1.36814029e-09-9.77801928e-14    2
 6.01459587e+04-1.09295466e+01-1.67820638e+00 4.25528459e-02-3.59188809e-05    3
 1.59603175e-08-2.88254684e-12 6.22946562e+04 3.08507210e+01                   4
C5H3                    C   5H   3          G    300.00   3500.00 1370.00      1
 1.06729929e+01 9.74586303e-03-3.33881731e-06 5.09387250e-10-2.86889364e-14    2
 6.39774214e+04-2.94129103e+01 3.35962353e+00 3.10987662e-02-2.67179083e-05    3
 1.18860739e-08-2.10472664e-12 6.59812846e+04 8.17219632e+00                   4
C5H2                    C   5H   2          G    300.00   3500.00 1260.00      1
 1.08586495e+01 8.25356564e-03-3.15379454e-06 5.51063165e-10-3.71272445e-14    2
 7.89908994e+04-3.35264725e+01 1.78531794e+00 3.70577928e-02-3.74445412e-05    3
 1.86943154e-08-3.63697887e-12 8.12773789e+04 1.23440607e+01                   4
C7H7O2                  C   7H   7O   2     G    300.00   3500.00 1420.00      1
 1.76964624e+01 2.58808959e-02-1.00755993e-05 1.78285133e-09-1.17592477e-13    2
 6.43630912e+03-6.45881470e+01-4.45172571e+00 8.82701582e-02-7.59797497e-05    3
 3.27237670e-08-5.56493678e-12 1.27263945e+04 5.00304722e+01                   4
O2C6H4CH3               C   7H   7O   2     G    300.00   3500.00 1300.00      1
 1.57011694e+01 2.91723897e-02-1.27991927e-05 2.73382155e-09-2.31734775e-13    2
 5.63564260e+03-5.46747931e+01-5.21645096e+00 9.35342985e-02-8.70629336e-05    3
 4.08177913e-08-7.55557510e-12 1.10742239e+04 5.17286697e+01                   4
OC6H4CH2                C   7H   6O   1     G    300.00   3500.00 1390.00      1
 1.45795344e+01 2.32519437e-02-8.58329374e-06 1.38947459e-09-7.81466978e-14    2
-5.01093183e+02-5.31869652e+01-4.82277789e+00 7.90859360e-02-6.88358034e-05    3
 3.02875607e-08-5.27564421e-12 4.89274964e+03 4.68072303e+01                   4
C6H5CH2O                C   7H   7O   1     G    300.00   3500.00 1650.00      1
 1.54569227e+01 2.51288522e-02-9.88344275e-06 1.85206220e-09-1.37473827e-13    2
 6.00712849e+03-5.64457004e+01-4.49397764e+00 7.34946712e-02-5.38523691e-05    3
 1.96172850e-08-2.82917425e-12 1.25909256e+04 4.97967788e+01                   4
BZCOOH                  C   7H   8O   2     G    300.00   3500.00 1550.00      1
 1.78036107e+01 3.06807111e-02-1.34555335e-05 2.81495359e-09-2.31878498e-13    2
-1.15055065e+04-6.47324084e+01-3.42659308e+00 8.54683337e-02-6.64758135e-05    3
 2.56193751e-08-3.91001099e-12-4.92414334e+03 4.69952939e+01                   4
C6H5O2                  C   6H   5O   2     G    300.00   3500.00 1300.00      1
 1.17436568e+01 2.50264983e-02-1.11158434e-05 2.39771212e-09-2.04780347e-13    2
 1.03023085e+04-3.29345583e+01-2.98072562e+00 7.03322902e-02-6.33917572e-05    3
 2.92058730e-08-5.36019591e-12 1.41306479e+04 4.19652270e+01                   4
C6H5CO                  C   7H   5O   1     G    300.00   3500.00 1470.00      1
 1.31799087e+01 2.42895707e-02-1.09067387e-05 2.35371847e-09-2.00195165e-13    2
 5.86598787e+03-4.37756649e+01-1.56203256e+00 6.44036967e-02-5.18395203e-05    3
 2.09173383e-08-3.35727336e-12 1.02001186e+04 3.30251959e+01                   4
RBBENZ                  C  14H  13          G    300.00   3500.00 1750.00      1
 5.34298872e+01-2.73976087e-03 1.40930517e-05-5.29858385e-09 5.98002535e-13    2
 9.33192272e+03-2.64139662e+02-8.67312060e+00 1.39209971e-01-1.07578147e-04    3
 4.10523491e-08-6.02355931e-12 3.10679755e+04 7.02252758e+01                   4
STILB                   C  14H  12          G    300.00   3500.00 1470.00      1
 3.31295358e+01 3.16424147e-02-7.88066874e-06 4.81370294e-10 4.43949926e-14    2
 1.37146851e+04-1.52659598e+02-1.11031623e+01 1.52003498e-01-1.30698101e-04    3
 5.61808860e-08-9.42831176e-12 2.67190984e+04 7.77787968e+01                   4
RBBENZOOH               C  14H  14O   2     G    300.00   3500.00 1390.00      1
 2.45960359e+01 6.70847362e-02-3.16552196e-05 7.12735227e-09-6.27188706e-13    2
-7.21416356e+03-9.76473229e+01-1.01910371e+01 1.67191421e-01-1.39684016e-04    3
 5.89397247e-08-9.94596073e-12 2.45664274e+03 8.16357090e+01                   4
RBBENZOO                C  14H  13O   2     G    300.00   3500.00 1370.00      1
 2.20515126e+01 6.70718760e-02-3.16675772e-05 7.13892279e-09-6.29044813e-13    2
 1.11280940e+04-8.22185224e+01-9.31390453e+00 1.58649736e-01-1.31935307e-04    3
 5.59310056e-08-9.53270956e-12 1.97222183e+04 7.89756546e+01                   4
QBBENZOOH               C  14H  13O   2     G    300.00   3500.00 1380.00      1
 2.50392782e+01 6.43939688e-02-3.06177262e-05 6.93819899e-09-6.13660452e-13    2
 1.02555756e+04-1.00870942e+02-8.15229194e+00 1.60601418e-01-1.35191041e-04    3
 5.74567086e-08-9.76556437e-12 1.94164490e+04 6.99496546e+01                   4
ZBBENZ                  C  14H  13O   4     G    300.00   3500.00 1360.00      1
 2.73944247e+01 6.88293330e-02-3.34701703e-05 7.71008172e-09-6.89822092e-13    2
-2.44016779e+03-1.05946545e+02-9.18072692e+00 1.76403308e-01-1.52117937e-04    3
 6.58707517e-08-1.13811217e-11 7.50827344e+03 8.17537182e+01                   4
KHYBBENZ                C  14H  12O   3     G    300.00   3500.00 1460.00      1
 2.68907577e+01 6.11068658e-02-2.84115712e-05 6.30145453e-09-5.47211887e-13    2
-2.19827626e+04-1.07049307e+02-7.41195553e+00 1.55086902e-01-1.24966403e-04    3
 5.03904188e-08-8.09669207e-12-1.19663704e+04 7.14228517e+01                   4
C14H13O                 C  14H  13O   1     G    300.00   3500.00 1450.00      1
 2.45301020e+01 5.83289648e-02-2.63012653e-05 5.70821145e-09-4.88285961e-13    2
 1.08230291e+04-9.99176314e+01-1.16317638e+01 1.58085836e-01-1.29498029e-04    3
 5.31549991e-08-8.66876660e-12 2.13099701e+04 8.79788989e+01                   4
C14H12O                 C  14H  12O   1     G    300.00   3500.00 1600.00      1
 2.85341713e+01 4.77197028e-02-1.97123161e-05 3.88726793e-09-3.03392983e-13    2
-1.40774973e+04-1.26522314e+02-8.99308371e+00 1.41537840e-01-1.07666820e-04    3
 4.05349779e-08-6.02959766e-12-2.06877575e+03 7.21629446e+01                   4
C5H5O                   C   5H   5O   1     G    300.00   3500.00 1450.00      1
 1.05801390e+01 2.13128784e-02-9.63052935e-06 2.09384798e-09-1.79321203e-13    2
 1.62543411e+04-3.26154734e+01-4.01979397e+00 6.15885556e-02-5.12950230e-05    3
 2.12499370e-08-3.48209517e-12 2.04883217e+04 4.32455666e+01                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459579e+00 2.39841575e-02-8.32755387e-06 8.47127652e-10 2.86249485e-14    2
 3.08659308e+03-9.73181555e+00-5.14379339e+00 6.04552343e-02-5.17455024e-05    3
 2.38195872e-08-4.52940274e-12 5.98166715e+03 4.83481227e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929577e+01 1.29021286e-02-2.02976642e-06-3.72417846e-10 8.59745728e-14    2
-2.22100459e+04-6.49015838e+01-5.23446578e+00 7.73770890e-02-7.06201498e-05    3
 3.20580235e-08-5.66410367e-12-1.58009124e+04 5.25540058e+01                   4
LC6H6                   C   6H   6          G    300.00   3500.00 1250.00      1
 1.28863876e+01 1.90072460e-02-7.30992558e-06 1.31482495e-09-9.21385787e-14    2
 3.55364843e+04-4.09021933e+01-1.05889383e+00 6.36321466e-02-6.08598062e-05    3
 2.98747613e-08-5.80412585e-12 3.90228046e+04 2.94875281e+01                   4
C6H4C2H3                C   8H   7          G    200.00   3500.00 1580.00      1
 1.99256075e+01 1.67315530e-02-4.18312961e-06 2.15370099e-10 3.07179808e-14    2
 3.89930312e+04-8.19571079e+01-3.96125911e+00 7.72046330e-02-6.15942816e-05    3
 2.44394849e-08-3.80221157e-12 4.65412811e+04 4.42096620e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155283e-02-1.38949871e-05 2.56768166e-09-1.71519559e-13    2
-2.17187243e+04-3.95715124e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733025e-12-1.73470426e+04 4.54334869e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353913e-06-2.12687588e-10 1.25840459e-13    2
-3.38086418e+03-4.22339552e+01-6.42956805e+00 9.31830717e-02-9.41722601e-05    3
 5.12938173e-08-1.10712258e-11 1.12339577e+03 5.49833260e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824814e+01 2.40796407e-02-4.51347945e-06-4.25076337e-10 1.44988489e-13    2
-3.97704754e+03-4.00543783e+01-6.60757189e+00 9.15233042e-02-9.24834753e-05    3
 5.05720227e-08-1.09413374e-11 4.82664709e+02 5.62014116e+01                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   3500.00 1450.00      1
 1.25818443e+01 2.64134519e-02-7.93799879e-06 4.38368240e-10 8.64078960e-14    2
-1.87828963e+04-3.81332333e+01-6.02884975e+00 7.77532977e-02-6.10481840e-05    3
 2.48568442e-08-4.12367417e-12-1.33857950e+04 5.85676633e+01                   4
C6H5C2H                 C   8H   6          G    200.00   3500.00 1280.00      1
 1.52608076e+01 2.33328927e-02-9.12947229e-06 1.67060897e-09-1.19620450e-13    2
 3.14643486e+04-5.61979008e+01-2.98097334e+00 8.03384582e-02-7.59328693e-05    3
 3.64640449e-08-6.91521341e-12 3.61342445e+04 3.63113150e+01                   4
C6H4C2H                 C   8H   5          G    200.00   3500.00 1410.00      1
 1.60102852e+01 1.80276839e-02-6.10631287e-06 8.89485624e-10-4.39310920e-14    2
 6.01004863e+04-5.91795508e+01-2.59308039e+00 7.08031891e-02-6.22504674e-05    3
 2.74351852e-08-4.75061541e-12 6.53466354e+04 3.69628594e+01                   4
C6H5C2H3                C   8H   8          G    200.00   3500.00 1620.00      1
 2.08689853e+01 1.76153525e-02-4.02709967e-06 7.62333198e-11 4.96213073e-14    2
 7.92336685e+03-8.97908225e+01-4.75261288e+00 8.08785579e-02-6.26041417e-05    3
 2.41820119e-08-3.67040626e-12 1.62247647e+04 4.61791070e+01                   4
C6H5C2H5                C   8H  10          G    200.00   3500.00 1660.00      1
 2.15526224e+01 2.25377527e-02-5.71678491e-06 3.25228910e-10 3.67333516e-14    2
-7.08672427e+03-9.37205827e+01-4.75947977e+00 8.59404087e-02-6.30083415e-05    3
 2.33338862e-08-3.42842587e-12 1.64889367e+03 4.65555372e+01                   4
C6H5C2H2                C   8H   7          G    200.00   3500.00 1520.00      1
 1.92541493e+01 1.80154928e-02-5.00513523e-06 4.35360010e-10 9.55509219e-15    2
 3.83998804e+04-7.81182474e+01-4.29898225e+00 7.99974179e-02-6.61715087e-05    3
 2.72627168e-08-4.40283911e-12 4.55600324e+04 4.53739369e+01                   4
C6H5CHCH3               C   8H   9          G    200.00   3500.00 1700.00      1
 2.17404159e+01 1.87953891e-02-4.10981050e-06 2.63146959e-14 6.24669644e-14    2
 1.18126541e+04-9.21825395e+01-3.04486857e+00 7.71137055e-02-5.55671485e-05    3
 2.01793745e-08-2.90508425e-12 2.02396509e+04 4.05439030e+01                   4
XYLENE                  C   8H  10          G    200.00   3500.00 1800.00      1
 2.00142025e+01 2.37296570e-02-6.76483884e-06 7.09529215e-10-1.05911394e-14    2
-8.30085767e+03-8.55893311e+01-3.92128796e+00 7.69196357e-02-5.10898211e-05    3
 1.71261893e-08-2.29068282e-12 3.15918887e+02 4.39545364e+01                   4
RXYLENE                 C   8H   9          G    200.00   3500.00 1620.00      1
 2.04972497e+01 2.14206934e-02-5.61362086e-06 3.90126528e-10 2.53125355e-14    2
 1.19614465e+04-8.71674754e+01-3.85447699e+00 8.15484138e-02-6.12874360e-05    3
 2.33011616e-08-3.51034102e-12 1.98514059e+04 4.20634392e+01                   4
INDENE                  C   9H   8          G    200.00   3500.00 1610.00      1
 2.31048443e+01 1.91297591e-02-4.53548120e-06 1.22196710e-10 5.15078704e-14    2
 8.53092089e+03-1.04304478e+02-6.87762290e+00 9.36203608e-02-7.39366630e-05    3
 2.88597461e-08-4.41084452e-12 1.81852753e+04 5.46222708e+01                   4
INDENYL                 C   9H   7          G    200.00   3500.00 1430.00      1
 2.02650248e+01 2.20602643e-02-7.28401475e-06 9.93375838e-10-4.12199482e-14    2
 2.49669757e+04-8.59379552e+01-6.82385337e+00 9.78333502e-02-8.67662727e-05    3
 3.80480416e-08-6.51930836e-12 3.27143949e+04 5.44392228e+01                   4
C10H7                   C  10H   7          G    200.00   3500.00 1490.00      1
 2.12397127e+01 2.27484190e-02-6.96640085e-06 8.04033892e-10-1.68765826e-14    2
 3.76445830e+04-9.11799918e+01-6.45168838e+00 9.70877508e-02-8.18046543e-05    3
 3.42887110e-08-5.63511100e-12 4.58966205e+04 5.34576808e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H7O                  C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C10H6CH3                C  11H   9          G    200.00   3500.00 1530.00      1
 2.52493034e+01 2.50352394e-02-6.91797176e-06 5.80757388e-10 1.70685087e-14    2
 3.22365770e+04-1.13732286e+02-6.94188403e+00 1.09195207e-01-8.94277435e-05    3
 3.65327276e-08-5.85743643e-12 4.20870803e+04 5.52614582e+01                   4
C10H7CH2                C  11H   9          G    200.00   3500.00 1480.00      1
 2.49658354e+01 2.73321443e-02-8.56500981e-06 1.05181516e-09-3.08784849e-14    2
 2.10853669e+04-1.11434350e+02-7.41870774e+00 1.14857936e-01-9.72735830e-05    3
 4.10106319e-08-6.78067861e-12 3.06711917e+04 5.74984546e+01                   4
C10H7CHO                C  11H   8O   1     G    200.00   3500.00 1700.00      1
 3.52801173e+01 1.31180999e-02-5.97608673e-07-9.89256296e-10 1.64132767e-13    2
-1.29136404e+04-1.70276910e+02-6.53399067e+00 1.11504236e-01-8.74089056e-05    3
 3.30543895e-08-4.84228574e-12 1.30315629e+03 5.36397371e+01                   4
C10H7CH3                C  11H  10          G    200.00   3500.00 1700.00      1
 3.19556671e+01 1.89589747e-02-2.92887930e-06-5.41537999e-10 1.30075116e-13    2
-1.51641167e+03-1.52538802e+02-7.17710534e+00 1.11036086e-01-8.41733896e-05    3
 3.13190543e-08-4.55530610e-12 1.17887310e+04 5.70191587e+01                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   3500.00 1800.00      1
 2.91191869e+01 2.86451308e-02-9.80098219e-06 1.51374083e-09-8.72237944e-14    2
-2.13626711e+04-1.32660114e+02-1.76841814e+00 9.72842531e-02-6.70002508e-05    3
 2.26986551e-08-3.02957300e-12-1.02431333e+04 3.45100483e+01                   4
CH3C10H6O               C  11H   9O   1     G    300.00   3500.00 1800.00      1
 2.60936624e+01 3.24954978e-02-1.30480618e-05 2.52260906e-09-1.95492396e-13    2
-2.87396993e+03-1.14905139e+02-1.85059487e+00 9.45938472e-02-6.47966864e-05    3
 2.16887663e-08-2.85745868e-12 7.18596268e+03 3.63350107e+01                   4
C12H8                   C  12H   8          G    200.00   3500.00 1570.00      1
 2.77000801e+01 2.26169409e-02-5.57154154e-06 2.34725133e-10 5.00956727e-14    2
 1.79557632e+04-1.32407942e+02-8.95027490e+00 1.15993641e-01-9.47849497e-05    3
 3.81172764e-08-5.98215771e-12 2.94639746e+04 6.09409166e+01                   4
C12H7                   C  12H   7          G    200.00   3500.00 1550.00      1
 2.72643903e+01 2.07706175e-02-5.09002112e-06 1.94274019e-10 4.95146521e-14    2
 5.03500896e+04-1.28964295e+02-8.21375630e+00 1.12327125e-01-9.36930927e-05    3
 3.83031220e-08-6.09707373e-12 6.13483151e+04 5.77457270e+01                   4
BIPHENYL                C  12H  10          G    200.00   3500.00 1620.00      1
 3.03550325e+01 2.42378629e-02-5.78855002e-06 1.73424746e-10 6.27217930e-14    2
 7.33500914e+03-1.42781766e+02-7.48580974e+00 1.17672041e-01-9.23016780e-05    3
 3.57755350e-08-5.43143103e-12 1.95954420e+04 5.80338349e+01                   4
C12H9                   C  12H   9          G    300.00   3500.00 1430.00      1
 2.37129726e+01 3.27032394e-02-1.16108739e-05 1.80515254e-09-1.00356247e-13    2
 4.00500330e+04-1.02303886e+02-9.58279779e+00 1.25838261e-01-1.09304953e-04    3
 4.73501777e-08-8.06277324e-12 4.95726233e+04 7.02380051e+01                   4
FLUORENE                C  13H  10          G    200.00   3500.00 1580.00      1
 3.04981916e+01 2.54134515e-02-6.12250971e-06 2.13473324e-10 6.26029969e-14    2
 6.42406071e+03-1.44876912e+02-9.12299946e+00 1.25720264e-01-1.01350497e-04    3
 4.03940585e-08-6.29508454e-12 1.89443571e+04 6.43961494e+01                   4
C6H5CH2C6H5             C  13H  12          G    200.00   3500.00 1730.00      1
 3.68978946e+01 2.09448951e-02-2.15140890e-06-1.01983322e-09 1.90993351e-13    2
 1.61235408e+03-1.77722051e+02-9.21937242e+00 1.27574414e-01-9.46047492e-05    3
 3.46076582e-08-4.95748807e-12 1.75689285e+04 7.00449656e+01                   4
C14H10                  C  14H  10          G    200.00   3500.00 1550.00      1
 3.33910328e+01 2.79675689e-02-7.16206046e-06 3.83005680e-10 5.29481034e-14    2
 8.53646106e+03-1.60739744e+02-9.79770356e+00 1.39422372e-01-1.15021548e-04    3
 4.67741830e-08-7.42949985e-12 2.19249693e+04 6.65486198e+01                   4
C14H9                   C  14H   9          G    298.15   3500.00 1380.00      1
 2.51054802e+01 4.12375730e-02-1.71094078e-05 3.35330065e-09-2.55891906e-13    2
 4.20489545e+04-1.12231128e+02-1.15966331e+01 1.47620510e-01-1.32743035e-04    3
 5.92149564e-08-1.03757571e-11 5.21787378e+04 7.66564976e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933977e+01 6.96117135e-02-3.71054121e-05 9.43826013e-09-9.32515879e-13    2
 4.61008358e+04-6.54256237e+01-1.33382684e+01 1.64875153e-01-1.52343443e-04    3
 7.13941909e-08-1.34236310e-11 5.34246890e+04 8.34001920e+01                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   3500.00 1170.00      1
 6.79293350e+00 9.36089894e-02-5.25184356e-05 1.38852184e-08-1.40951794e-12    2
 1.04787082e+04-8.65156268e+00-1.16088786e+01 1.56521167e-01-1.33175074e-04    3
 5.98434170e-08-1.12296458e-11 1.47847322e+04 8.30156967e+01                   4
C16H10                  C  16H  10          G    200.00   3500.00 1560.00      1
 3.81807346e+01 2.83119223e-02-6.73305412e-06 1.57165250e-10 8.21178663e-14    2
 9.09208909e+03-1.88517714e+02-1.17161985e+01 1.56252776e-01-1.29753106e-04    3
 5.27298370e-08-8.34298979e-12 2.46599322e+04 7.43946040e+01                   4
BENZYNE                 C   6H   4          G    300.00   3500.00 1400.00      1
 1.09465819e+01 1.50373246e-02-5.27844959e-06 8.14607580e-10-4.49073365e-14    2
 5.03301418e+04-3.53782934e+01-3.73796173e+00 5.69931634e-02-5.02311341e-05    3
 2.22206478e-08-3.86741452e-12 5.44418140e+04 4.04070822e+01                   4
LC6H5                   C   6H   5          G    300.00   3500.00 1140.00      1
 1.23076076e+01 1.68261952e-02-6.51181370e-06 1.21158891e-09-8.99428216e-14    2
 5.89425072e+04-3.55373249e+01 1.67614173e-01 5.94226632e-02-6.25597980e-05    3
 3.39881879e-08-7.27779348e-12 6.17104257e+04 2.46218079e+01                   4
C6H2                    C   6H   2          G    200.00   3500.00  700.00      1
 9.95239962e+00 1.43744770e-02-7.32585544e-06 1.80931771e-09-1.74471744e-13    2
 8.06473020e+04-2.49945457e+01-5.39476473e-01 7.43280546e-02-1.35797808e-04    3
 1.24163558e-07-4.38724146e-11 8.21161647e+04 2.18805022e+01                   4
C6H3                    C   6H   3          G    300.00   3500.00 1320.00      1
 1.19194523e+01 1.16137832e-02-4.19264522e-06 6.84693072e-10-4.17887567e-14    2
 8.26280760e+04-3.29876543e+01 4.46601450e+00 3.41999583e-02-2.98587533e-05    3
 1.36473739e-08-2.49684195e-12 8.45957836e+04 5.04018537e+00                   4
C6H4                    C   6H   4          G    300.00   3500.00 1360.00      1
 1.74447675e+01 6.21306707e-03-9.80963855e-07 8.00594627e-11-2.88320761e-15    2
 5.49568894e+04-6.59208082e+01-1.17305610e+00 6.09713718e-02-6.13761529e-05    3
 2.96855443e-08-5.44506791e-12 6.00209374e+04 2.96241244e+01                   4
C8H2                    C   8H   2          G    300.00   3500.00 1060.00      1
 1.62719352e+01 9.99874490e-03-2.93037079e-06 2.89537337e-10 2.52406325e-16    2
 1.07885460e+05-5.89733614e+01 1.87361717e-01 7.06952485e-02-8.88216494e-05    3
 5.43092094e-08-1.27402363e-11 1.11295389e+05 1.95626382e+01                   4
BIN1B                   C  20H  10          G    300.00   3500.00 1780.00      1
-5.70256700e+00 1.43432300e-01-8.80724700e-05 2.76799200e-08-3.52289900e-12    2
 2.77808900e+04 4.34481200e+01-5.70256700e+00 1.43432300e-01-8.80724700e-05    3
 2.76799200e-08-3.52289900e-12 2.77808900e+04 4.34481200e+01                   4
BIN1A                   C  20H  16          G    300.00   3500.00 1780.00      1
-3.24173600e+00 1.58222900e-01-9.46183500e-05 2.81843100e-08-3.56131000e-12    2
 2.17869900e+04 3.00825300e+01-3.24173600e+00 1.58222900e-01-9.46183500e-05    3
 2.81843100e-08-3.56131000e-12 2.17869900e+04 3.00825300e+01                   4
RMCYC6                  C   7H  13          G    300.00   3500.00 1800.00      1
 1.73339062e+01 3.85260822e-02-1.58310821e-05 3.15191459e-09-2.53163787e-13    2
-5.89957980e+03-7.33836420e+01-9.95790329e+00 9.91745477e-02-6.63714701e-05    3
 2.18705768e-08-2.85297798e-12 3.92547162e+03 7.43253244e+01                   4
MCYC6                   C   7H  14          G    300.00   3500.00 1800.00      1
 1.67194568e+01 4.36180644e-02-1.87773363e-05 3.92059022e-09-3.26702983e-13    2
-2.91866300e+04-7.40611878e+01-1.01006358e+01 1.03218270e-01-6.84441744e-05    3
 2.23157154e-08-2.88158149e-12-1.95313967e+04 7.10947481e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623566e-02-8.52218598e-06 1.36123710e-09-7.97159889e-14    2
-5.90596972e+03-6.59480381e+01-8.70136947e+00 9.66875823e-02-8.77887356e-05    3
 3.96542563e-08-7.01685714e-12 1.03797027e+03 6.35339364e+01                   4
RC9H11                  C   9H  11          G    300.00   3500.00 1800.00      1
 1.94777671e+01 3.52558917e-02-1.42493230e-05 2.76058348e-09-2.13045169e-13    2
 6.10938819e+03-7.94713741e+01-1.83523003e+00 8.26181075e-02-5.37178363e-05    3
 1.73785513e-08-2.24331848e-12 1.37820672e+04 3.58790126e+01                   4
TMBENZ                  C   9H  12          G    300.00   3500.00 1800.00      1
 1.47576861e+01 4.50315825e-02-1.97554195e-05 4.21197817e-09-3.57314917e-13    2
-1.09025839e+04-5.35378398e+01-2.75522789e+00 8.39491691e-02-5.21867417e-05    3
 1.62235790e-08-2.02559281e-12-4.59793488e+03 4.12457040e+01                   4
NPBENZ                  C   9H  12          G    300.00   3500.00 1600.00      1
 1.88963371e+01 3.80090295e-02-1.52789389e-05 2.95630099e-09-2.27699217e-13    2
-8.96605283e+03-7.62711275e+01-5.58650157e+00 9.92161261e-02-7.26605920e-05    3
 2.68653231e-08-3.96348393e-12-1.13154446e+03 5.33514397e+01                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934216e-02-1.83631832e-05 3.88491135e-09-3.27420808e-13    2
 4.39687821e+03-8.23923218e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836943e-12 1.50954180e+04 7.84485932e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565535e-05 2.20632462e-09-1.51941205e-13    2
-9.85314331e+03-1.11161770e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
DCYC5                   C  10H  16          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748171e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
ODECAL                  C  10H  18          G    300.00   3500.00 1800.00      1
 2.82109941e+01 4.74108396e-02-1.82963852e-05 3.42084161e-09-2.57817125e-13    2
-2.68355230e+04-1.31410203e+02-1.02710769e+01 1.32926553e-01-8.95594797e-05    3
 2.98145803e-08-3.92361417e-12-1.29819774e+04 7.68627930e+01                   4
DECALIN                 C  10H  18          G    300.00   3500.00 1750.00      1
 2.70110296e+01 4.68748171e-02-1.63895490e-05 2.62563687e-09-1.59789734e-13    2
-3.79226289e+04-1.35167747e+02-1.45870783e+01 1.41956207e-01-9.78878828e-05    3
 3.36726212e-08-4.59507321e-12-2.33632912e+04 8.87980358e+01                   4
NC10H20                 C  10H  20          G    300.00   3500.00 1800.00      1
 2.82971791e+01 4.89478938e-02-1.82737062e-05 3.23575201e-09-2.26811843e-13    2
-3.12534582e+04-1.16784058e+02-2.31417710e+00 1.16973130e-01-7.49614029e-05    3
 2.42311952e-08-3.14284562e-12-2.02333700e+04 4.88909878e+01                   4
NC10MOOH                C  10H  20O   2     G    300.00   3500.00 1790.00      1
 2.73219585e+01 3.55870996e-02-1.24650774e-05 2.00089264e-09-1.21997682e-13    2
-4.84634178e+04-1.12262056e+02 1.16215154e+00 9.40447688e-02-6.14519510e-05    3
 2.02455383e-08-2.67013255e-12-3.90982069e+04 2.91745387e+01                   4
NC10H22                 C  10H  22          G    300.00   3500.00 1800.00      1
 2.92878918e+01 5.29920990e-02-1.98404553e-05 3.55616370e-09-2.54281184e-13    2
-4.56232379e+04-1.22752047e+02-2.17870143e+00 1.22917862e-01-7.81119243e-05    3
 2.51381893e-08-3.25178473e-12-3.42952643e+04 4.75517200e+01                   4
DIBZFUR                 C  12H   8O   1     G    300.00   3500.00 1410.00      1
 2.49525256e+01 3.24730728e-02-1.15459374e-05 1.79679054e-09-9.97833661e-14    2
-5.30753651e+03-1.13355893e+02-1.16970901e+01 1.36443614e-01-1.22152896e-04    3
 5.40932248e-08-9.37220078e-12 5.02765510e+03 7.60497478e+01                   4
NC12H26                 C  12H  26          G    300.00   3500.00 1800.00      1
 3.61414095e+01 6.11045883e-02-2.24641073e-05 3.93182440e-09-2.73349362e-13    2
-5.40359186e+04-1.56831960e+02-2.66627705e+00 1.47343892e-01-9.43301934e-05    3
 3.05488933e-08-3.97016449e-12-4.00651514e+04 5.32033350e+01                   4
IC16H34                 C  16H  34          G    300.00   3500.00 1590.00      1
 4.72524600e+01 8.54680758e-02-3.36612723e-05 6.38202029e-09-4.82094887e-13    2
-7.78744143e+04-2.24182950e+02-9.93612249e+00 2.29338723e-01-1.69388298e-04    3
 6.32906266e-08-9.42998896e-12-5.96884450e+04 7.82391931e+01                   4
NC16H34                 C  16H  34          G    300.00   3500.00 1800.00      1
 4.98210237e+01 7.73881687e-02-2.77557896e-05 4.69678103e-09-3.12959242e-13    2
-7.08514664e+04-2.24842855e+02-3.64057977e+00 1.96191732e-01-1.26758759e-04    3
 4.13645475e-08-5.40570458e-12-5.16052891e+04 6.45024955e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835937e-02-9.17249481e-06 1.42952536e-09-8.46466182e-14    2
 3.95646504e+03-1.44540610e+02-1.09331575e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619032e+01-7.89283135e-03 1.09697207e-05-3.89489830e-09 4.38586294e-13    2
-1.76924159e+04-2.71823424e+02-1.36343924e+01 1.41210048e-01-1.13282679e-04    3
 4.21245088e-08-5.95299803e-12 6.46225047e+03 9.13157248e+01                   4
RDECALIN                C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620334e+01 4.11366392e-02-1.36024110e-05 2.01592782e-09-1.09376625e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278109e+00 9.04971362e+01                   4
RODECA                  C  10H  17          G    300.00   3500.00 1800.00      1
 2.85620334e+01 4.11366392e-02-1.36024110e-05 2.01592782e-09-1.09376625e-13    2
-1.53025063e+04-1.39641687e+02-1.39601308e+01 1.35630337e-01-9.23471594e-05    3
 3.11806495e-08-4.16003241e-12 5.47278109e+00 9.04971362e+01                   4
NC10H19                 C  10H  19          G    300.00   3500.00 1800.00      1
 9.88287390e+00 2.86275350e-02-1.23662428e-05 2.58308509e-09-2.14520963e-13    2
 7.14211639e+03-2.81379758e+01-9.61360662e-01 5.27258341e-02-3.24481586e-05    3
 1.00208317e-08-1.24754133e-12 1.10460408e+04 3.05532839e+01                   4
NC10H21                 C  10H  21          G    300.00   3500.00 1800.00      1
 2.63212692e+01 5.52219738e-02-2.21266526e-05 4.33498891e-09-3.42316503e-13    2
-2.10175171e+04-1.03192977e+02-1.81057271e+00 1.17737178e-01-7.42226562e-05    3
 2.36298050e-08-3.02215208e-12-1.08900540e+04 4.90624204e+01                   4
NC12H25                 C  12H  25          G    300.00   3500.00 1800.00      1
 3.17005579e+01 6.61544325e-02-2.66295230e-05 5.21804509e-09-4.10998518e-13    2
-2.88525898e+04-1.31607624e+02-2.06085145e+00 1.41179787e-01-8.91506513e-05    3
 2.83740186e-08-3.62710595e-12-1.66984825e+04 5.11161660e+01                   4
IC16H33                 C  16H  33          G    300.00   3500.00 1650.00      1
 5.11453588e+01 7.53296743e-02-2.79263242e-05 4.92908201e-09-3.44364401e-13    2
-5.61938874e+04-2.43048234e+02-8.95216175e+00 2.21020633e-01-1.60372651e-04    3
 5.84427492e-08-8.45249580e-12-3.63617056e+04 7.69829165e+01                   4
NC16H33                 C  16H  33          G    300.00   3500.00 1800.00      1
 4.66278372e+01 8.00212238e-02-3.03236334e-05 5.55903616e-09-4.09822553e-13    2
-4.61545210e+04-2.04019480e+02-3.22413374e+00 1.90803381e-01-1.22642098e-04    3
 3.97510601e-08-5.15871477e-12-2.82078115e+04 6.57897858e+01                   4
BIN1C                   C  20H   4          G   300.00   4000.00  1000.00      1
 .279698426e+02 .447047097e-01-.165223093e-04 .275199987e-08-.171198257e-12    2
-.832698077e+04-.148330566e+03-.841721188e+01 .122499448e+00-.329768495e-04    3
-.527684334e-07 .303949355e-10 .241443283e+04 .443201113e+02                   4
BIN2A                   C  40H  31          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .397395323e+03-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .283409758e+05 .136281912e+03                   4
BIN2B                   C  40H  16          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
-.435148944e+04-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .195176885e+05 .109755604e+03                   4
BIN2C                   C  40H   8          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
-.170085815e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .447424565e+04 .886402226e+02                   4
BIN3A                   C  80H  60          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .303189596e+04-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .578481001e+05 .254746237e+03                   4
BIN3B                   C  80H  24          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
-.213600710e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .239919342e+05 .198395827e+03                   4
BIN3C                   C  80H   8          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
-.466742552e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09-.609495158e+04 .156165064e+03                   4
BIN4A                   C 160H 116          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .105380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .118028497e+06 .473857298e+03                   4
BIN4B                   C 160H  32          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.680343262e+05-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .178969826e+05 .354560890e+03                   4
BIN4C                   C 160H   8          G   300.00   4000.00  1000.00      1
 .203770010e+03 .325689326e+00-.120370758e-03 .200492744e-07-.124723874e-11    2
-.106005602e+06-.113404212e+04-.651786613e+02 .882711219e+00-.164645194e-03    3
-.476244713e-06 .251238312e-09-.272333461e+05 .291214746e+03                   4
BIN5A                   C 320H 224          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .352119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .247380465e+06 .927804457e+03                   4
BIN5B                   C 320H  64          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.135714032e+06-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .361485852e+05 .709121781e+03                   4
BIN5C                   C 320H  16          G   300.00   4000.00  1000.00      1
 .407540019e+03 .651378652e+00-.240741515e-03 .400985487e-07-.249447749e-11    2
-.212011205e+06-.226808424e+04-.130357323e+03 .176542244e+01-.329290388e-03    3
-.952489427e-06 .502476624e-09-.544666921e+05 .582429491e+03                   4
BIN6A                   C 640H 432          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .909146192e+05-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .507419557e+06 .173874832e+04                   4
BIN6B                   C 640H 128          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.271428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .722971705e+05 .141824356e+04                   4
BIN6C                   C 640H  32          G   300.00   4000.00  1000.00      1
 .815080039e+03 .130275730e+01-.481483031e-03 .801970974e-07-.498895498e-11    2
-.424022410e+06-.453616849e+04-.260714645e+03 .353084488e+01-.658580775e-03    3
-.190497885e-05 .100495325e-08-.108933384e+06 .116485898e+04                   4
BIN7A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          813
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .219703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .101891965e+07 .319868647e+04                   4
BIN7B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          250
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.528501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .142639667e+06 .276398698e+04                   4
BIN7C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           63
 .159241877e+04 .254519198e+01-.940671563e-03 .156680764e-06-.974690233e-11    2
-.826135381e+06-.886271923e+04-.509037242e+03 .689863702e+01-.129017531e-02    3
-.371755916e-05 .196193239e-08-.210676521e+06 .227342492e+04                   4
BIN8A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1563
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .525439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .209454960e+07 .599019956e+04                   4
BIN8B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          500
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.106037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .282300003e+06 .554001391e+04                   4
BIN8C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          125
 .318395553e+04 .508897425e+01-.188082211e-02 .313274746e-06-.194884061e-10    2
-.165482925e+07-.177213274e+05-.101820055e+04 .137927917e+02-.257439985e-02    3
-.743934801e-05 .392490001e-08-.424111287e+06 .454722041e+04                   4
BIN9A                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         3000
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .105415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .433609933e+07 .163588732e+05                   4
BIN9B                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         1000
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.212075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .564600007e+06 .110800278e+05                   4
BIN9C                   C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          250
 .636791107e+04 .101779485e+02-.376164423e-02 .626549492e-06-.389768122e-10    2
-.330965851e+07-.354426549e+05-.203640111e+04 .275855833e+02-.514879970e-02    3
-.148786960e-04 .784980002e-08-.848222575e+06 .909444082e+04                   4
BIN10A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5750
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .171313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .820225091e+07 .320518708e+05                   4
BIN10B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         2000
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.424150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .112920001e+07 .221600556e+05                   4
BIN10C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          500
 .127356256e+05 .203555829e+02-.752317236e-02 .125307965e-05-.779524215e-10    2
-.662269050e+07-.708776326e+05-.407366633e+04 .551694512e+02-.102903246e-01    3
-.297652946e-04 .157023945e-07-.169942448e+07 .182009216e+05                   4
BIN11A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        11000
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .262917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .154586477e+08 .627960702e+05                   4
BIN11B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         4000
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.848301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .225840003e+07 .443201113e+05                   4
BIN11C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         1000
 .254712512e+05 .407111657e+02-.150463447e-01 .250615929e-05-.155904843e-09    2
-.132453810e+08-.141755265e+06-.814733266e+04 .110338902e+03-.205806492e-01    3
-.595305892e-04 .314047890e-07-.339884896e+07 .364018432e+05                   4
BIN12A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        21000
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .367089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290315457e+08 .122952718e+06                   4
BIN12B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         8000
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169660271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .451680005e+07 .886402226e+05                   4
BIN12C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         2000
 .509425024e+05 .814223315e+02-.300926894e-01 .501231859e-05-.311809686e-09    2
-.264907620e+08-.283510531e+06-.162946653e+05 .220677805e+03-.411612984e-01    3
-.119061178e-03 .628095780e-07-.679769791e+07 .728036864e+05                   4
BIN13A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        40000
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .416688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .542915920e+08 .240626590e+06                   4
BIN13B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        16000
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.339320543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .903360011e+07 .177280445e+06                   4
BIN13C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         4000
 .101885005e+06 .162844663e+03-.601853789e-01 .100246372e-04-.623619372e-09    2
-.529815240e+08-.567021061e+06-.325893306e+05 .441355610e+03-.823225969e-01    3
-.238122357e-03 .125619156e-06-.135953958e+08 .145607373e+06                   4
BIN14A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        76000
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .198394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101040185e+09 .470695489e+06                   4
BIN14B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        32000
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678641086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .180672002e+08 .354560890e+06                   4
BIN14C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         8000
 .203770010e+06 .325689326e+03-.120370758e+00 .200492744e-04-.124723874e-08    2
-.105963048e+09-.113404212e+07-.651786613e+05 .882711219e+03-.164645194e+00    3
-.476244713e-03 .251238312e-06-.271907917e+08 .291214746e+06                   4
BIN15A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       144000
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.873175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .186994373e+09 .920275597e+06                   4
BIN15B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        64000
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135728217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361344004e+08 .709121781e+06                   4
BIN15C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        16000
 .407540019e+06 .651378652e+03-.240741515e+00 .400985487e-04-.249447749e-08    2
-.211926096e+09-.226808424e+07-.130357323e+06 .176542244e+04-.329290388e+00    3
-.952489427e-03 .502476624e-06-.543815833e+08 .582429491e+06                   4
BIN16A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       272000
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428627973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343816752e+09 .179832043e+07                   4
BIN16B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       128000
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271456434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .722688009e+08 .141824356e+07                   4
BIN16C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        32000
 .815080039e+06 .130275730e+04-.481483031e+00 .801970974e-04-.498895498e-08    2
-.423852192e+09-.453616849e+07-.260714645e+06 .353084488e+04-.658580775e+00    3
-.190497885e-02 .100495325e-05-.108763167e+09 .116485898e+07                   4
BIN17A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       500000
 .195633111e+07 .312683969e+04-.115564137e+01 .192486706e-03-.119743423e-07    2
-.133324395e+09-.981860207e+07-.548565677e+06 .866959432e+04-.309406979e+01    3
-.273451411e-02 .181552901e-05 .612587417e+09 .342986263e+07                   4
BIN17B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       250000
 .174811516e+07 .279404436e+04-.103264433e+01 .171999992e-03-.106998911e-07    2
-.530188348e+09-.927066036e+07-.526075742e+06 .765621551e+04-.206105310e+01    3
-.329802709e-02 .189968347e-05 .141150002e+09 .277000696e+07                   4
BIN17C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H        62500
 .159195320e+07 .254444786e+04-.940396545e+00 .156634956e-03-.974405269e-08    2
-.827836313e+09-.885970408e+07-.509208291e+06 .689618140e+04-.128629058e+01    3
-.372066182e-02 .196279931e-05-.212428060e+09 .227511520e+07                   4
BIN18A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       937500
 .386060824e+07 .617048055e+04-.228053348e+01 .379851734e-03-.236300717e-07    2
-.365864779e+09-.195002187e+08-.109150887e+07 .170858439e+05-.592988540e+01    3
-.560990646e-02 .365209663e-05 .110731548e+10 .669476134e+07                   4
BIN18B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       500000
 .349623033e+07 .558808872e+04-.206528866e+01 .343999983e-03-.213997822e-07    2
-.106037670e+10-.185413207e+08-.105215148e+07 .153124310e+05-.412210619e+01    3
-.659605418e-02 .379936694e-05 .282300003e+09 .554001391e+07                   4
BIN18C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       125000
 .318390640e+07 .508889572e+04-.188079309e+01 .313269912e-03-.194881054e-07    2
-.165567263e+10-.177194082e+08-.101841658e+07 .137923628e+05-.257258115e+01    3
-.744132365e-02 .392559863e-05-.424856120e+09 .455023040e+07                   4
BIN19A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1750000
 .761710851e+07 .121745634e+05-.449956845e+01 .749460110e-03-.466229179e-07    2
-.930161534e+09-.387264666e+08-.217177277e+07 .336649985e+05-.113432625e+02    3
-.115015694e-01 .734627050e-05 .197891225e+10 .130595948e+08                   4
BIN19B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1000000
 .699246065e+07 .111761774e+05-.413057731e+01 .687999967e-03-.427995643e-07    2
-.212075339e+10-.370826415e+08-.210430297e+07 .306248620e+05-.824421238e+01    3
-.131921084e-01 .759873388e-05 .564600007e+09 .110800278e+08                   4
BIN19C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       250000
 .636781280e+07 .101777914e+05-.376158618e+01 .626539824e-03-.389762108e-07    2
-.331134525e+10-.354388163e+08-.203683317e+07 .275847256e+05-.514516230e+01    3
-.148826473e-01 .785119726e-05-.849712239e+09 .910046080e+07                   4
BIN20A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      3250000
 .150260011e+08 .240163315e+05-.887613985e+01 .147843351e-02-.919713846e-07    2
-.225718702e+10-.769049915e+08-.432105561e+07 .663166181e+05-.216535082e+02    3
-.235666518e-01 .147766955e-04 .348638709e+10 .254593340e+08                   4
BIN20B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      2000000
 .139849213e+08 .223523549e+05-.826115463e+01 .137599993e-02-.855991287e-07    2
-.424150678e+10-.741652829e+08-.420860594e+07 .612497241e+05-.164884248e+02    3
-.263842167e-01 .151974678e-04 .112920001e+10 .221600556e+08                   4
BIN20C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H       500000
 .127356256e+08 .203555829e+05-.752317236e+01 .125307965e-02-.779524215e-07    2
-.662269050e+10-.708776326e+08-.407366633e+07 .551694512e+05-.102903246e+02    3
-.297652946e-01 .157023945e-04-.169942448e+10 .182009216e+08                   4
BIN21A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      6000000
 .296355702e+08 .473670724e+05-.175062856e+02 .291589358e-02-.181393867e-06    2
-.530810195e+10-.152714099e+09-.859713135e+07 .130606479e+06-.412409831e+02    3
-.482603296e-01 .297216998e-04 .602989935e+10 .495989567e+08                   4
BIN21B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      4000000
 .279698426e+08 .447047097e+05-.165223093e+02 .275199987e-02-.171198257e-06    2
-.848301357e+10-.148330566e+09-.841721188e+07 .122499448e+06-.329768495e+02    3
-.527684334e-01 .303949355e-04 .225840003e+10 .443201113e+08                   4
BIN21C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      1000000
 .254712512e+08 .407111657e+05-.150463447e+02 .250615929e-02-.155904843e-06    2
-.132453810e+11-.141755265e+09-.814733266e+07 .110338902e+06-.205806492e+02    3
-.595305892e-01 .314047890e-04-.339884896e+10 .364018432e+08                   4
BIN22A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H     12000000
 .592711404e+08 .947341447e+05-.350125712e+02 .583178717e-02-.362787734e-06    2
-.106162039e+11-.305428199e+09-.171942627e+08 .261212957e+06-.824819661e+02    3
-.965206591e-01 .594433996e-04 .120597987e+11 .991979134e+08                   4
BIN22B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      8000000
 .559396852e+08 .894094194e+05-.330446185e+02 .550399973e-02-.342396515e-06    2
-.169660271e+11-.296661132e+09-.168344238e+08 .244998896e+06-.659536990e+02    3
-.105536867e+00 .607898710e-04 .451680005e+10 .886402226e+08                   4
BIN22C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      2000000
 .509425024e+08 .814223315e+05-.300926894e+02 .501231859e-02-.311809686e-06    2
-.264907620e+11-.283510531e+09-.162946653e+08 .220677805e+06-.411612984e+02    3
-.119061178e+00 .628095780e-04-.679769791e+10 .728036864e+08                   4
BIN23A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     24000000
 .118542281e+09 .189468289e+06-.700251424e+02 .116635743e-01-.725575467e-06    2
-.212324078e+11-.610856398e+09-.343885254e+08 .522425915e+06-.164963932e+03    3
-.193041318e+00 .118886799e-03 .241195974e+11 .198395827e+09                   4
BIN23B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     16000000
 .111879370e+09 .178818839e+06-.660892370e+02 .110079995e-01-.684793029e-06    2
-.339320543e+11-.593322263e+09-.336688475e+08 .489997793e+06-.131907398e+03    3
-.211073734e+00 .121579742e-03 .903360011e+10 .177280445e+09                   4
BIN23C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H      4000000
 .101885005e+09 .162844663e+06-.601853789e+02 .100246372e-01-.623619372e-06    2
-.529815240e+11-.567021061e+09-.325893306e+08 .441355610e+06-.823225969e+02    3
-.238122357e+00 .125619156e-03-.135953958e+11 .145607373e+09                   4
BIN24A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     48000000
 .237084562e+09 .378936579e+06-.140050285e+03 .233271487e-01-.145115093e-05    2
-.424648156e+11-.122171280e+10-.687770508e+08 .104485183e+07-.329927864e+03    3
-.386082637e+00 .237773599e-03 .482391948e+11 .396791654e+09                   4
BIN24B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     32000000
 .223758741e+09 .357637678e+06-.132178474e+03 .220159989e-01-.136958606e-05    2
-.678641086e+11-.118664453e+10-.673376950e+08 .979995585e+06-.263814796e+03    3
-.422147467e+00 .243159484e-03 .180672002e+11 .354560890e+09                   4
BIN24C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H      8000000
 .203770010e+09 .325689326e+06-.120370758e+03 .200492744e-01-.124723874e-05    2
-.105963048e+12-.113404212e+10-.651786613e+08 .882711219e+06-.164645194e+03    3
-.476244713e+00 .251238312e-03-.271907917e+11 .291214746e+09                   4
BIN25A                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     96000000
 .474169124e+09 .757873158e+06-.280100570e+03 .466542973e-01-.290230187e-05    2
-.849296311e+11-.244342559e+10-.137554102e+09 .208970366e+07-.659855729e+03    3
-.772165273e+00 .475547197e-03 .964783896e+11 .793583307e+09                   4
BIN25B                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     64000000
 .447517482e+09 .715275356e+06-.264356948e+03 .440319979e-01-.273917212e-05    2
-.135728217e+12-.237328905e+10-.134675390e+09 .195999117e+07-.527629592e+03    3
-.844294935e+00 .486318968e-03 .361344004e+11 .709121781e+09                   4
BIN25C                  C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     16000000
 .407540019e+09 .651378652e+06-.240741515e+03 .400985487e-01-.249447749e-05    2
-.211926096e+12-.226808424e+10-.130357323e+09 .176542244e+07-.329290388e+03    3
-.952489427e+00 .502476624e-03-.543815833e+11 .582429491e+09                   4
BIN1AJ                  C  20H  15          G   300.00   4000.00  1000.00      1
 .384004130e+02 .613760802e-01-.226838420e-04 .377828116e-08-.235041851e-12    2
 .583425289e+05-.190858878e+03-.946290891e+01 .179252381e+00-.989756752e-04    3
-.116559979e-07 .214782048e-10 .722142317e+05 .597553003e+02                   4
BIN1BJ                  C  20H   9          G   300.00   4000.00  1000.00      1
 .329670254e+02 .526917977e-01-.194742383e-04 .324368101e-08-.201785086e-12    2
 .610771833e+05-.161481167e+03-.895697031e+01 .146820540e+00-.577692501e-04    3
-.392441219e-07 .283752285e-10 .736083600e+05 .601566475e+02                   4
BIN1CJ                  C  20H   3          G   300.00   4000.00  1000.00      1
 .279698426e+02 .447047097e-01-.165223093e-04 .275199987e-08-.171198257e-12    2
 .516730192e+05-.148330566e+03-.841721188e+01 .122499448e+00-.329768495e-04    3
-.527684334e-07 .303949355e-10 .624144328e+05 .443201113e+02                   4
BIN2AJ                  C  40H  30          G   300.00   4000.00  1000.00      1
 .759883346e+02 .121453540e+00-.448877300e-04 .747661988e-08-.465110589e-12    2
 .603973953e+05-.376351286e+03-.224069955e+02 .373191638e+00-.228373343e-03    3
 .179614865e-08 .353583380e-10 .883409758e+05 .136281912e+03                   4
BIN2BJ                  C  40H  15          G   300.00   4000.00  1000.00      1
 .626025956e+02 .100058870e+00-.369805239e-04 .615957460e-08-.383178953e-12    2
 .556485106e+05-.314195266e+03-.175541017e+02 .277427018e+00-.990102332e-04    3
-.875044514e-07 .580969283e-10 .795176885e+05 .109755604e+03                   4
BIN2CJ                  C  40H   7          G   300.00   4000.00  1000.00      1
 .559396852e+02 .894094194e-01-.330446185e-04 .550399973e-08-.342396515e-12    2
 .429914185e+05-.296661132e+03-.168344238e+02 .244998896e+00-.659536990e-04    3
-.105536867e-06 .607898710e-10 .644742457e+05 .886402226e+02                   4
BIN3AJ                  C  80H  59          G   300.00   4000.00  1000.00      1
 .150797478e+03 .241022357e+00-.890788896e-04 .148372172e-07-.923003567e-12    2
 .630318960e+05-.764406699e+03-.455633619e+02 .756332498e+00-.489114578e-03    3
 .351844886e-07 .598168799e-10 .117848100e+06 .254746237e+03                   4
BIN3BJ                  C  80H  23          G   300.00   4000.00  1000.00      1
 .118542281e+03 .189468289e+00-.700251424e-04 .116635743e-07-.725575467e-12    2
 .386399290e+05-.610856398e+03-.343885254e+02 .522425915e+00-.164963932e-03    3
-.193041318e-06 .118886799e-09 .839919342e+05 .198395827e+03                   4
BIN3CJ                  C  80H   7          G   300.00   4000.00  1000.00      1
 .105216460e+03 .168169388e+00-.621533316e-04 .103524246e-07-.644010591e-12    2
 .133257448e+05-.575788129e+03-.329491696e+02 .457569671e+00-.988508639e-04    3
-.229106149e-06 .124272685e-09 .539050484e+05 .156165064e+03                   4
BIN4AJ                  C 160H 115          G   300.00   4000.00  1000.00      1
 .299236573e+03 .478275269e+00-.176764639e-03 .294423892e-07-.183157191e-11    2
 .705380025e+05-.155222165e+04-.926254655e+02 .153256344e+01-.104296494e-02    3
 .133553360e-06 .978341677e-10 .178028497e+06 .473857298e+03                   4
BIN4BJ                  C 160H  31          G   300.00   4000.00  1000.00      1
 .223758741e+03 .357637678e+00-.132178474e-03 .220159989e-07-.136958606e-11    2
-.803432616e+04-.118664453e+04-.673376950e+02 .979995585e+00-.263814796e-03    3
-.422147467e-06 .243159484e-09 .778969826e+05 .354560890e+03                   4
BIN4CJ                  C 160H   7          G   300.00   4000.00  1000.00      1
 .203770010e+03 .325689326e+00-.120370758e-03 .200492744e-07-.124723874e-11    2
-.460056024e+05-.113404212e+04-.651786613e+02 .882711219e+00-.164645194e-03    3
-.476244713e-06 .251238312e-09 .327666539e+05 .291214746e+03                   4
BIN5AJ                  C 320H 223          G   300.00   4000.00  1000.00      1
 .593310588e+03 .948299129e+00-.350479658e-03 .583768256e-07-.363154476e-11    2
 .952119959e+05-.312882274e+04-.194461399e+03 .312434830e+01-.224387754e-02    3
 .412099583e-06 .147772804e-09 .307380465e+06 .927804457e+03                   4
BIN5BJ                  C 320H  63          G   300.00   4000.00  1000.00      1
 .447517482e+03 .715275356e+00-.264356948e-03 .440319979e-07-.273917212e-11    2
-.757140323e+05-.237328905e+04-.134675390e+03 .195999117e+01-.527629592e-03    3
-.844294935e-06 .486318968e-09 .961485852e+05 .709121781e+03                   4
BIN5CJ                  C 320H  15          G   300.00   4000.00  1000.00      1
 .407540019e+03 .651378652e+00-.240741515e-03 .400985487e-07-.249447749e-11    2
-.152011205e+06-.226808424e+04-.130357323e+03 .176542244e+01-.329290388e-03    3
-.952489427e-06 .502476624e-09 .553330788e+04 .582429491e+03                   4
BIN6AJ                  C 640H 431          G   300.00   4000.00  1000.00      1
 .117696475e+04 .188116422e+01-.695255086e-03 .115803539e-06-.720398434e-11    2
 .150914619e+06-.634005997e+04-.398024258e+03 .633800264e+01-.476093625e-02    3
 .108624875e-05 .206199066e-09 .567419557e+06 .173874832e+04                   4
BIN6BJ                  C 640H 127          G   300.00   4000.00  1000.00      1
 .895034964e+03 .143055071e+01-.528713896e-03 .880639958e-07-.547834423e-11    2
-.211428065e+06-.474657811e+04-.269350780e+03 .391998234e+01-.105525918e-02    3
-.168858987e-05 .972637936e-09 .132297170e+06 .141824356e+04                   4
BIN6CJ                  C 640H  31          G   300.00   4000.00  1000.00      1
 .815080039e+03 .130275730e+01-.481483031e-03 .801970974e-07-.498895498e-11    2
-.364022410e+06-.453616849e+04-.260714645e+03 .353084488e+01-.658580775e-03    3
-.190497885e-05 .100495325e-08-.489333842e+05 .116485898e+04                   4
BIN7AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          812
 .227996401e+04 .364410804e+01-.134681737e-02 .224329490e-06-.139552395e-10    2
 .279703936e+06-.125294003e+05-.798183644e+03 .125608657e+02-.983885162e-02    3
 .263510017e-05 .228737231e-09 .107891965e+07 .319868647e+04                   4
BIN7BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H          249
 .174821343e+04 .279420142e+01-.103270238e-02 .172009660e-06-.107004925e-10    2
-.468501603e+06-.927449889e+04-.525643684e+03 .765707323e+01-.206469049e-02    3
-.329407582e-05 .189828623e-08 .202639667e+06 .276398698e+04                   4
BIN7CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         1250 H           62
 .159241877e+04 .254519198e+01-.940671563e-03 .156680764e-06-.974690233e-11    2
-.766135381e+06-.886271923e+04-.509037242e+03 .689863702e+01-.129017531e-02    3
-.371755916e-05 .196193239e-08-.150676521e+06 .227342492e+04                   4
BIN8AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H         1562
 .452144611e+04 .722670975e+01-.267090277e-02 .444872681e-06-.276749385e-10    2
 .585439399e+06-.253601694e+05-.163861142e+04 .254934056e+02-.207827201e-01    3
 .632122666e-05 .101241844e-09 .215454960e+07 .599019956e+04                   4
BIN8BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          499
 .349623033e+04 .558808872e+01-.206528866e-02 .343999983e-06-.213997822e-10    2
-.100037670e+07-.185413207e+05-.105215148e+04 .153124310e+02-.412210619e-02    3
-.659605418e-05 .379936694e-08 .342300003e+06 .554001391e+04                   4
BIN8CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         2500 H          124
 .318395553e+04 .508897425e+01-.188082211e-02 .313274746e-06-.194884061e-10    2
-.159482925e+07-.177213274e+05-.101820055e+04 .137927917e+02-.257439985e-02    3
-.743934801e-05 .392490001e-08-.364111287e+06 .454722041e+04                   4
BIN9AJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H         2999
 .865818826e+04 .138385401e+02-.511455367e-02 .851893682e-06-.529951738e-10    2
 .111415823e+07-.414661751e+05-.228422245e+04 .387318925e+02-.165083459e-01    3
-.868400451e-05 .692549819e-08 .439609933e+07 .163588732e+05                   4
BIN9BJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          999
 .699246065e+04 .111761774e+02-.413057731e-02 .687999967e-06-.427995643e-10    2
-.206075339e+07-.370826415e+05-.210430297e+04 .306248620e+02-.824421238e-02    3
-.131921084e-04 .759873388e-08 .624600007e+06 .110800278e+05                   4
BIN9CJ                  C   0H   0          G   300.00   4000.00  1000.00      1&
C         5000 H          249
 .636791107e+04 .101779485e+02-.376164423e-02 .626549492e-06-.389768122e-10    2
-.324965851e+07-.354426549e+05-.203640111e+04 .275855833e+02-.514879970e-02    3
-.148786960e-04 .784980002e-08-.788222575e+06 .909444082e+04                   4
BIN10AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         5749
 .171082588e+05 .273444419e+02-.101061683e-01 .168331032e-05-.104716498e-09    2
 .177313926e+07-.823882471e+05-.454552290e+04 .764512640e+02-.319873125e-01    3
-.179275707e-04 .139337536e-07 .826225091e+07 .320518708e+05                   4
BIN10BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H         1999
 .139849213e+05 .223523549e+02-.826115463e-02 .137599993e-05-.855991287e-10    2
-.418150678e+07-.741652829e+05-.420860594e+04 .612497241e+02-.164884248e-01    3
-.263842167e-04 .151974678e-07 .118920001e+07 .221600556e+05                   4
BIN10CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        10000 H          499
 .127356256e+05 .203555829e+02-.752317236e-02 .125307965e-05-.779524215e-10    2
-.656269050e+07-.708776326e+05-.407366633e+04 .551694512e+02-.102903246e-01    3
-.297652946e-04 .157023945e-07-.163942448e+07 .182009216e+05                   4
BIN11AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H        10999
 .337998892e+05 .540229790e+02-.199662265e-01 .332562787e-05-.206882891e-09    2
 .268917711e+07-.163672934e+06-.904693005e+04 .150874055e+03-.619013169e-01    3
-.369900700e-04 .280386106e-07 .155186477e+08 .627960702e+05                   4
BIN11BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H         3999
 .279698426e+05 .447047097e+02-.165223093e-01 .275199987e-05-.171198257e-09    2
-.842301357e+07-.148330566e+06-.841721188e+04 .122499448e+03-.329768495e-01    3
-.527684334e-04 .303949355e-07 .231840003e+07 .443201113e+05                   4
BIN11CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        20000 H          999
 .254712512e+05 .407111657e+02-.150463447e-01 .250615929e-05-.155904843e-09    2
-.131853810e+08-.141755265e+06-.814733266e+04 .110338902e+03-.205806492e-01    3
-.595305892e-04 .314047890e-07-.333884896e+07 .364018432e+05                   4
BIN12AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H        20999
 .667669147e+05 .106714777e+03-.394404648e-01 .656930888e-05-.408667976e-09    2
 .373089841e+07-.325154101e+06-.180039004e+05 .297694595e+03-.119670567e+00    3
-.762341918e-04 .564138391e-07 .290915457e+08 .122952718e+06                   4
BIN12BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         7999
 .559396852e+05 .894094194e+02-.330446185e-01 .550399973e-05-.342396515e-09    2
-.169060271e+08-.296661132e+06-.168344238e+05 .244998896e+03-.659536990e-01    3
-.105536867e-03 .607898710e-07 .457680005e+07 .886402226e+05                   4
BIN12CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        40000 H         1999
 .509425024e+05 .814223315e+02-.300926894e-01 .501231859e-05-.311809686e-09    2
-.264307620e+08-.283510531e+06-.162946653e+05 .220677805e+03-.411612984e-01    3
-.119061178e-03 .628095780e-07-.673769791e+07 .728036864e+05                   4
BIN13AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        39999
 .131868102e+06 .210767191e+03-.778969533e-01 .129747241e-04-.807140343e-09    2
 .422688521e+07-.645924667e+06-.358278812e+05 .587282159e+03-.231077001e+00    3
-.156976488e-03 .113500914e-06 .543515920e+08 .240626590e+06                   4
BIN13BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H        15999
 .111879370e+06 .178818839e+03-.660892370e-01 .110079995e-04-.684793029e-09    2
-.338720543e+08-.593322263e+06-.336688475e+05 .489997793e+03-.131907398e+00    3
-.211073734e-03 .121579742e-06 .909360011e+07 .177280445e+06                   4
BIN13CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C        80000 H         3999
 .101885005e+06 .162844663e+03-.601853789e-01 .100246372e-04-.623619372e-09    2
-.529215240e+08-.567021061e+06-.325893306e+05 .441355610e+03-.823225969e-01    3
-.238122357e-03 .125619156e-06-.135353958e+08 .145607373e+06                   4
BIN14AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        75999
 .260404748e+06 .416209656e+03-.153825954e+00 .256216607e-04-.159388947e-08    2
 .204394716e+07-.128308227e+07-.712959235e+05 .115835026e+04-.445625734e+00    3
-.322969183e-03 .228348299e-06 .101100185e+09 .470695489e+06                   4
BIN14BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H        31999
 .223758741e+06 .357637678e+03-.132178474e+00 .220159989e-04-.136958606e-08    2
-.678041086e+08-.118664453e+07-.673376950e+05 .979995585e+03-.263814796e+00    3
-.422147467e-03 .243159484e-06 .181272002e+08 .354560890e+06                   4
BIN14CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       160000 H         7999
 .203770010e+06 .325689326e+03-.120370758e+00 .200492744e-04-.124723874e-08    2
-.105903048e+09-.113404212e+07-.651786613e+05 .882711219e+03-.164645194e+00    3
-.476244713e-03 .251238312e-06-.271307917e+08 .291214746e+06                   4
BIN15AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H       143999
 .514146586e+06 .821769862e+03-.303716002e+00 .505877465e-04-.314699650e-08    2
-.867175217e+07-.254863040e+07-.141872169e+06 .228427239e+04-.858194934e+00    3
-.663970781e-03 .459389541e-06 .187054373e+09 .920275597e+06                   4
BIN15BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        63999
 .447517482e+06 .715275356e+03-.264356948e+00 .440319979e-04-.273917212e-08    2
-.135668217e+09-.237328905e+07-.134675390e+06 .195999117e+04-.527629592e+00    3
-.844294935e-03 .486318968e-06 .361944004e+08 .709121781e+06                   4
BIN15CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       320000 H        15999
 .407540019e+06 .651378652e+03-.240741515e+00 .400985487e-04-.249447749e-08    2
-.211866096e+09-.226808424e+07-.130357323e+06 .176542244e+04-.329290388e+00    3
-.952489427e-03 .502476624e-06-.543215833e+08 .582429491e+06                   4
BIN16AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       271999
 .101496735e+07 .162224082e+04-.599560194e+00 .998643433e-04-.621242812e-08    2
-.428027973e+08-.506219253e+07-.282304982e+06 .450368854e+04-.165027680e+01    3
-.136400639e-02 .924164967e-06 .343876752e+09 .179832043e+07                   4
BIN16BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H       127999
 .895034964e+06 .143055071e+04-.528713896e+00 .880639958e-04-.547834423e-08    2
-.271396434e+09-.474657811e+07-.269350780e+06 .391998234e+04-.105525918e+01    3
-.168858987e-02 .972637936e-06 .723288009e+08 .141824356e+07                   4
BIN16CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C       640000 H        31999
 .815080039e+06 .130275730e+04-.481483031e+00 .801970974e-04-.498895498e-08    2
-.423792192e+09-.453616849e+07-.260714645e+06 .353084488e+04-.658580775e+00    3
-.190497885e-02 .100495325e-05-.108703167e+09 .116485898e+07                   4
BIN17AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       499999
 .195633111e+07 .312683969e+04-.115564137e+01 .192486706e-03-.119743423e-07    2
-.133264395e+09-.981860207e+07-.548565677e+06 .866959432e+04-.309406979e+01    3
-.273451411e-02 .181552901e-05 .612647417e+09 .342986263e+07                   4
BIN17BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H       249999
 .174811516e+07 .279404436e+04-.103264433e+01 .171999992e-03-.106998911e-07    2
-.530128348e+09-.927066036e+07-.526075742e+06 .765621551e+04-.206105310e+01    3
-.329802709e-02 .189968347e-05 .141210002e+09 .277000696e+07                   4
BIN17CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      1250000 H        62499
 .159195320e+07 .254444786e+04-.940396545e+00 .156634956e-03-.974405269e-08    2
-.827776313e+09-.885970408e+07-.509208291e+06 .689618140e+04-.128629058e+01    3
-.372066182e-02 .196279931e-05-.212368060e+09 .227511520e+07                   4
BIN18AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       937499
 .386060824e+07 .617048055e+04-.228053348e+01 .379851734e-03-.236300717e-07    2
-.365804779e+09-.195002187e+08-.109150887e+07 .170858439e+05-.592988540e+01    3
-.560990646e-02 .365209663e-05 .110737548e+10 .669476134e+07                   4
BIN18BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       499999
 .349623033e+07 .558808872e+04-.206528866e+01 .343999983e-03-.213997822e-07    2
-.106031670e+10-.185413207e+08-.105215148e+07 .153124310e+05-.412210619e+01    3
-.659605418e-02 .379936694e-05 .282360003e+09 .554001391e+07                   4
BIN18CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      2500000 H       124999
 .318390640e+07 .508889572e+04-.188079309e+01 .313269912e-03-.194881054e-07    2
-.165561263e+10-.177194082e+08-.101841658e+07 .137923628e+05-.257258115e+01    3
-.744132365e-02 .392559863e-05-.424796120e+09 .455023040e+07                   4
BIN19AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H      1749999
 .761710851e+07 .121745634e+05-.449956845e+01 .749460110e-03-.466229179e-07    2
-.930101534e+09-.387264666e+08-.217177277e+07 .336649985e+05-.113432625e+02    3
-.115015694e-01 .734627050e-05 .197897225e+10 .130595948e+08                   4
BIN19BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       999999
 .699246065e+07 .111761774e+05-.413057731e+01 .687999967e-03-.427995643e-07    2
-.212069339e+10-.370826415e+08-.210430297e+07 .306248620e+05-.824421238e+01    3
-.131921084e-01 .759873388e-05 .564660007e+09 .110800278e+08                   4
BIN19CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C      5000000 H       249999
 .636781280e+07 .101777914e+05-.376158618e+01 .626539824e-03-.389762108e-07    2
-.331128525e+10-.354388163e+08-.203683317e+07 .275847256e+05-.514516230e+01    3
-.148826473e-01 .785119726e-05-.849652239e+09 .910046080e+07                   4
BIN20AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      3249999
 .150260011e+08 .240163315e+05-.887613985e+01 .147843351e-02-.919713846e-07    2
-.225712702e+10-.769049915e+08-.432105561e+07 .663166181e+05-.216535082e+02    3
-.235666518e-01 .147766955e-04 .348644709e+10 .254593340e+08                   4
BIN20BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H      1999999
 .139849213e+08 .223523549e+05-.826115463e+01 .137599993e-02-.855991287e-07    2
-.424144678e+10-.741652829e+08-.420860594e+07 .612497241e+05-.164884248e+02    3
-.263842167e-01 .151974678e-04 .112926001e+10 .221600556e+08                   4
BIN20CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     10000000 H       499999
 .127356256e+08 .203555829e+05-.752317236e+01 .125307965e-02-.779524215e-07    2
-.662263050e+10-.708776326e+08-.407366633e+07 .551694512e+05-.102903246e+02    3
-.297652946e-01 .157023945e-04-.169936448e+10 .182009216e+08                   4
BIN21AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      5999999
 .296355702e+08 .473670724e+05-.175062856e+02 .291589358e-02-.181393867e-06    2
-.530804195e+10-.152714099e+09-.859713135e+07 .130606479e+06-.412409831e+02    3
-.482603296e-01 .297216998e-04 .602995935e+10 .495989567e+08                   4
BIN21BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H      3999999
 .279698426e+08 .447047097e+05-.165223093e+02 .275199987e-02-.171198257e-06    2
-.848295357e+10-.148330566e+09-.841721188e+07 .122499448e+06-.329768495e+02    3
-.527684334e-01 .303949355e-04 .225846003e+10 .443201113e+08                   4
BIN21CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     20000000 H       999999
 .254712512e+08 .407111657e+05-.150463447e+02 .250615929e-02-.155904843e-06    2
-.132453210e+11-.141755265e+09-.814733266e+07 .110338902e+06-.205806492e+02    3
-.595305892e-01 .314047890e-04-.339878896e+10 .364018432e+08                   4
BIN22AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H     11999999
 .592711404e+08 .947341447e+05-.350125712e+02 .583178717e-02-.362787734e-06    2
-.106161439e+11-.305428199e+09-.171942627e+08 .261212957e+06-.824819661e+02    3
-.965206591e-01 .594433996e-04 .120598587e+11 .991979134e+08                   4
BIN22BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      7999999
 .559396852e+08 .894094194e+05-.330446185e+02 .550399973e-02-.342396515e-06    2
-.169659671e+11-.296661132e+09-.168344238e+08 .244998896e+06-.659536990e+02    3
-.105536867e+00 .607898710e-04 .451686005e+10 .886402226e+08                   4
BIN22CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     40000000 H      1999999
 .509425024e+08 .814223315e+05-.300926894e+02 .501231859e-02-.311809686e-06    2
-.264907020e+11-.283510531e+09-.162946653e+08 .220677805e+06-.411612984e+02    3
-.119061178e+00 .628095780e-04-.679763791e+10 .728036864e+08                   4
BIN23AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     23999999
 .118542281e+09 .189468289e+06-.700251424e+02 .116635743e-01-.725575467e-06    2
-.212323478e+11-.610856398e+09-.343885254e+08 .522425915e+06-.164963932e+03    3
-.193041318e+00 .118886799e-03 .241196574e+11 .198395827e+09                   4
BIN23BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H     15999999
 .111879370e+09 .178818839e+06-.660892370e+02 .110079995e-01-.684793029e-06    2
-.339319943e+11-.593322263e+09-.336688475e+08 .489997793e+06-.131907398e+03    3
-.211073734e+00 .121579742e-03 .903366011e+10 .177280445e+09                   4
BIN23CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C     80000000 H      3999999
 .101885005e+09 .162844663e+06-.601853789e+02 .100246372e-01-.623619372e-06    2
-.529814640e+11-.567021061e+09-.325893306e+08 .441355610e+06-.823225969e+02    3
-.238122357e+00 .125619156e-03-.135953358e+11 .145607373e+09                   4
BIN24AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     47999999
 .237084562e+09 .378936579e+06-.140050285e+03 .233271487e-01-.145115093e-05    2
-.424647556e+11-.122171280e+10-.687770508e+08 .104485183e+07-.329927864e+03    3
-.386082637e+00 .237773599e-03 .482392548e+11 .396791654e+09                   4
BIN24BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H     31999999
 .223758741e+09 .357637678e+06-.132178474e+03 .220159989e-01-.136958606e-05    2
-.678640486e+11-.118664453e+10-.673376950e+08 .979995585e+06-.263814796e+03    3
-.422147467e+00 .243159484e-03 .180672602e+11 .354560890e+09                   4
BIN24CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    160000000 H      7999999
 .203770010e+09 .325689326e+06-.120370758e+03 .200492744e-01-.124723874e-05    2
-.105962988e+12-.113404212e+10-.651786613e+08 .882711219e+06-.164645194e+03    3
-.476244713e+00 .251238312e-03-.271907317e+11 .291214746e+09                   4
BIN25AJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     95999999
 .474169124e+09 .757873158e+06-.280100570e+03 .466542973e-01-.290230187e-05    2
-.849295711e+11-.244342559e+10-.137554102e+09 .208970366e+07-.659855729e+03    3
-.772165273e+00 .475547197e-03 .964784496e+11 .793583307e+09                   4
BIN25BJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     63999999
 .447517482e+09 .715275356e+06-.264356948e+03 .440319979e-01-.273917212e-05    2
-.135728157e+12-.237328905e+10-.134675390e+09 .195999117e+07-.527629592e+03    3
-.844294935e+00 .486318968e-03 .361344604e+11 .709121781e+09                   4
BIN25CJ                 C   0H   0          G   300.00   4000.00  1000.00      1&
C    320000000 H     15999999
 .407540019e+09 .651378652e+06-.240741515e+03 .400985487e-01-.249447749e-05    2
-.211926036e+12-.226808424e+10-.130357323e+09 .176542244e+07-.329290388e+03    3
-.952489427e+00 .502476624e-03-.543815233e+11 .582429491e+09                   4
CSOLID                  C   1               G    300.00   4000.00 1000.00      1
 .159828070E+01 .143065097E-02-.509435105E-06 .864401302E-10-.534349530E-14    2
-.745940284E+03-.930332005E+01-.303744539E+00 .436036227E-02 .198268825E-05    3
-.643472598E-08 .299601320E-11-.109458288E+03 .108301475E+01                   4
END
