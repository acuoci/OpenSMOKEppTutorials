!***********************************************************************
!SURFACE MECHANISM OF POX of CH4 on PT wire gauze
!***********************************************************************      
!****                                                                  *     
!****     CH4-O2 SURFACE MECHANISM  ON PT                              *    
!****                                                                  *         
!****     Version 1.0   Spring 2005                                    *
!****                                                                  *         
!****     Raul Quiceno, Olaf Deutschmann, IWR, Heidelberg University,  *
!****     Germany            *                                         *
!****     Contact: mail@detchem.com (O. Deutschmann)                   *
!****                                                                  *
!****     Reference:                                                   *
!****     R. Quiceno, J. Perez-Ramyrez, J. Warnatz, O. Deutschmann.    *
!****     Appl. Catal. A: General (2006)                               *
!****     www.detchem.com/mechanisms                                   *
!****                                                                  *
!****                                                                  *
!****     Kinetic data format: DETCHEM                                 *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****      STICK: A in next reaction is initial sticking coefficient   *
!****                                                                  *
!****      $..  : additional coverage dependence of Ea (3rd column)    *
!****               or changed reaction order (2nd column)             *
!****                                                                  *
!****      see manuals on www.detchem.com for details                  *
!****                                                                  *
!****      The kinetic data of the backward reactions of               *
!****      reactions in Section 3 are calculated                       *
!****      from thermodynamics (k_b = k_f /K)                          *
!****                                                                  *
!****     Surface site density: 2.72E-9 mol/cm**2                      *
!****                                                                  *
!****     CHEMKIN format                                               *
!****                                                                  *
!***********************************************************************

THERMO
   300.000  1000.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2            (adjust)  N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
C2H3O             T 9/92C   2H   3O   1    0G   298.150  3500.000 1000.00      1
 0.48131470E+00 0.20711914E-01-0.12693155E-04 0.34579642E-08-0.35399703E-12    2
 0.15648642E+05 0.34629876E+02 0.10854772E+01 0.12845259E-01 0.24138660E-05    3
-0.44642672E-08-0.29381916E-12 0.15910655E+05 0.33395312E+02 0.16817588E+05    4
C2H4              121286C   2H   4          G  0300.00   5000.00  1000.00      1
 0.03528418E+02 0.11485185E-01-0.04418385E-04 0.07844600E-08-0.05266848E-12    2
 0.04428288E+05 0.02230389E+02-0.08614880E+01 0.02796162E+00-0.03388677E-03    3
 0.02785152E-06-0.09737879E-10 0.05573046E+05 0.02421148E+03                   4
C2H5               12387C   2H   5          G  0300.00   5000.00  1000.00      1
 0.07190480E+02 0.06484077E-01-0.06428064E-05-0.02347879E-08 0.03880877E-12    2
 0.10674549E+05-0.14780892E+02 0.02690701E+02 0.08719133E-01 0.04419838E-04    3
 0.09338703E-08-0.03927773E-10 0.12870404E+05 0.12138195E+02                   4
C2H5O2             MAR97C   2H   5O   2    0G   300.000  5000.000 1401.00      1
 1.01174925E+01 1.14414478E-02-3.87093107E-06 5.96456991E-10-3.44195189E-14    2
-6.72193488E+03-2.51029911E+01 1.14509259E+00 3.40950493E-02-2.63317159E-05    3
 1.09211311E-08-1.86974412E-12-3.75862702E+03 2.25106527E+01                   4
C2H5OOH                 C   2H   6O   2    0G   300.000  5000.000 1409.000     1
 1.26555265E+01 1.13347220E-02-3.82256729E-06 5.88089793E-10-3.39112055E-14    2
-2.63839689E+04-4.04200223E+01 1.76442089E-01 4.29475359E-02-3.45056187E-05    3
 1.40909800E-08-2.29710196E-12-2.23628129E+04 2.56156874E+01                   4
C2H6              121686C   2H   6          G  0300.00   4000.00  1000.00      1
 0.04825938E+02 0.13840429E-01-0.04557258E-04 0.06724967E-08-0.03598161E-12    2
-0.12717793E+05-0.05239506E+02 0.14625388E+01 0.15494667E-01 0.05780507E-04    3
-0.12578319E-07 0.04586267E-10-0.11239176E+05 0.14432295E+02                   4
CH2O              121286C   1H   2O   1     G  0300.00   5000.00  1000.00      1
 0.02995606E+02 0.06681321E-01-0.02628954E-04 0.04737153E-08-0.03212517E-12    2
-0.15320369E+05 0.06912572E+02 0.16527311E+01 0.12631439E-01-0.01888168E-03    3
 0.02050031E-06-0.08413237E-10-0.14865404E+05 0.13784820E+02                   4
CH2OH              MAR97C   1H   3O   1     G   300.00   5000.00  1410.00      1
 6.00127803E+00 4.98721568E-03-1.60953515E-06 2.40227135E-10-1.35582700E-14    2
-3.50157098E+03-6.92836844E+00 2.60067849E+00 1.28447854E-02-8.33796185E-06    3
 2.75727606E-09-3.57041106E-13-2.33478724E+03 1.13272307E+01                   4
CH3               121286C   1H   3          G  0300.00   5000.00  1000.00      1
 0.02844051E+02 0.06137974E-01-0.02230345E-04 0.03785161E-08-0.02452159E-12    2
 0.16437809E+05 0.05452697E+02 0.02430442E+02 0.11124099E-01-0.01680220E-03    3
 0.16218288E-07-0.05864952E-10 0.16423781E+05 0.06789794E+02                   4
CH3CHO     9/20/ 1      C   2H   4O   1    0G   300.000  5000.000 1366.000     1
 7.06734034E+00 9.72785577E-03-3.36197228E-06 5.25639518E-10-3.06473991E-14    2
-2.32754287E+04-1.33686458E+01 1.98023941E+00 1.69300955E-02-4.36472545E-06    3
-1.70119601E-09 7.72360943E-13-2.10195065E+04 1.56487028E+01                   4
CH3CO             120186C   2H   3O   1     G  0300.00   5000.00  1000.00      1
 0.05612279E+02 0.08449886E-01-0.02854147E-04 0.04238376E-08-0.02268404E-12    2
-0.05187863E+05-0.03274949E+02 0.03125278E+02 0.09778220E-01 0.04521448E-04    3
-0.09009462E-07 0.03193718E-10-0.04108508E+05 0.01122885E+03                   4
CH3O              121686C   1H   3O   1     G  0300.00   3000.00  1000.00      1
 0.03770799E+02 0.07871497E-01-0.02656384E-04 0.03944431E-08-0.02112616E-12    2
 0.12783252E+03 0.02929575E+02 0.02106204E+02 0.07216595E-01 0.05338472E-04    3
-0.07377636E-07 0.02075610E-10 0.09786011E+04 0.13152177E+02                   4
CH3O2             BURCT C   1H   3O   2    0G   300.000  5000.000 1000.00      1
 0.66812963E+01 0.80057271E-02-0.27188507E-05 0.40631365E-09-0.21927725E-13    2
 0.52621851E+03-0.99423847E+01 0.20986490E+01 0.15786357E-01 0.75683261E-07    3
-0.11274587E-07 0.56665133E-11 0.20695879E+04 0.15007068E+02                   4
CH3O2H  CH4O2     T 5/92C   1H   4O   2    0G   298.150  5000.000 1000.00      1
 0.66499943E+01 0.10351461E-01-0.33524105E-05 0.53645535E-09-0.33949756E-13    2
-0.19232344E+05-0.77922626E+01 0.27586279E+01 0.18150526E-01-0.40892298E-05    3
-0.68391987E-08 0.41430701E-11-0.17986394E+05 0.13071986E+02-0.16404863E+05    4
CH3OH             121686C   1H   4O   1     G  0300.00   5000.00  1000.00      1
 0.04029061E+02 0.09376593E-01-0.03050254E-04 0.04358793E-08-0.02224723E-12    2
-0.02615791E+06 0.02378196E+02 0.02660115E+02 0.07341508E-01 0.07170051E-04    3
-0.08793194E-07 0.02390570E-10-0.02535348E+06 0.01123263E+03                   4
CH4                     C   1H   4    0    0G  0300.00   5000.00  1000.00      1
 1.68347883E+00 1.02372356E-02-3.87512864E-06 6.78558487E-10-4.50342312E-14    2
-1.00807871E+04 9.62339497E+00 7.78741479E-01 1.74766835E-02-2.78340904E-05    3
 3.04970804E-08-1.22393068E-11-9.82522852E+03 1.37221947E+01                   4
CHO      HCO      121286H   1C   1O   1     G  0300.00   5000.00  1000.00      1
 0.03557271E+02 0.03345572E-01-0.13350060E-05 0.02470572E-08-0.01713850E-12    2
 0.03916324E+05 0.05552299E+02 0.02898329E+02 0.06199146E-01-0.09623084E-04    3
 0.10898249E-07-0.04574885E-10 0.04159922E+05 0.08983614E+02                   4
CO                      C   1O   1    0    0G  0300.00   5000.00  1000.00      1
 3.02507806E+00 1.44268852E-03-5.63082779E-07 1.01858133E-10-6.91095156E-15    2
-1.42683496E+04 6.10821772E+00 3.26245165E+00 1.51194085E-03-3.88175522E-06    3
 5.58194424E-09-2.47495123E-12-1.43105391E+04 4.84889698E+00                   4
CO2                     C   1O   2    0    0G  0300.00   5000.00  1000.00      1
 4.45362282E+00 3.14016873E-03-1.27841054E-06 2.39399667E-10-1.66903319E-14    2
-4.89669609E+04-9.55395877E-01 2.27572465E+00 9.92207229E-03-1.04091132E-05    3
 6.86668678E-09-2.11728009E-12-4.83731406E+04 1.01884880E+01                   4
DC2OOH1           T10/10C  2 H  5 O  2    0 G   200.000  6000.000  1000.00     1
 8.88872432E+00 1.35833179E-02-4.91116949E-06 7.92343362E-10-4.73525704E-14    2
-7.44107388E+03-1.90789836E+01 4.50099327E+00 6.87965342E-03 4.74143971E-05    3
-6.92287127E-08 2.87395324E-11-5.39547911E+03 7.91490068E+00-3.45206633E+03    4
H                 120186H   1               G  0300.00   5000.00  1000.00      1
 0.02500000E+02 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.02547162E+06-0.04601176E+01 0.02500000E+02 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.02547162E+06-0.04601176E+01                   4
H2                121286H   2               G  0300.00   5000.00  1000.00      1
 0.02991423E+02 0.07000644E-02-0.05633828E-06-0.09231578E-10 0.15827519E-14    2
-0.08350340E+04-0.13551101E+01 0.03298124E+02 0.08249441E-02-0.08143015E-05    3
-0.09475434E-09 0.04134872E-11-0.10125209E+04-0.03294094E+02                   4
H2O                20387H   2O   1          G  0300.00   5000.00  1000.00      1
 0.02672145E+02 0.03056293E-01-0.08730260E-05 0.12009964E-09-0.06391618E-13    2
-0.02989921E+06 0.06862817E+02 0.03386842E+02 0.03474982E-01-0.06354696E-04    3
 0.06968581E-07-0.02506588E-10-0.03020811E+06 0.02590232E+02                   4
H2O2              120186H   2O   2          G  0300.00   5000.00  1000.00      1
 0.04573167E+02 0.04336136E-01-0.14746888E-05 0.02348903E-08-0.14316536E-13    2
-0.01800696E+06 0.05011369E+01 0.03388753E+02 0.06569226E-01-0.14850125E-06    3
-0.04625805E-07 0.02471514E-10-0.01766314E+06 0.06785363E+02                   4
HO2                20387H   1O   2          G  0300.00   5000.00  1000.00      1
 0.04072191E+02 0.02131296E-01-0.05308145E-05 0.06112269E-09-0.02841164E-13    2
-0.15797270E+03 0.03476029E+02 0.02979963E+02 0.04996697E-01-0.03790997E-04    3
 0.02354192E-07-0.08089024E-11 0.01762273E+04 0.09222724E+02                   4
O                 120186O   1               G  0300.00   5000.00  1000.00      1
 0.02542059E+02-0.02755061E-03-0.03102803E-07 0.04551067E-10-0.04368051E-14    2
 0.02923080E+06 0.04920308E+02 0.02946428E+02-0.16381665E-02 0.02421031E-04    3
-0.16028431E-08 0.03890696E-11 0.02914764E+06 0.02963995E+02                   4
O2                121386O   2               G  0300.00   5000.00  1000.00      1
 0.03697578E+02 0.06135197E-02-0.12588420E-06 0.01775281E-09-0.11364354E-14    2
-0.12339301E+04 0.03189165E+02 0.03212936E+02 0.11274864E-02-0.05756150E-05    3
 0.13138773E-08-0.08768554E-11-0.10052490E+04 0.06034737E+02                   4
OH                121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 0.03886888E+05 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 0.03606781E+05 0.13588605E+01                   4
OXIRAN            L 8/88C   2H   4O   1    0G   200.000  6000.000 1000.00      1
 0.54887641E+01 0.12046190E-01-0.43336931E-05 0.70028311E-09-0.41949088E-13    2
-0.91804251E+04-0.70799605E+01 0.37590532E+01-0.94412180E-02 0.80309721E-04    3
-0.10080788E-06 0.40039921E-10-0.75608143E+04 0.78497475E+01-0.63304657E+04    4
C_Pt                   0C   1PT  1          I    300.00   3000.00 1000.00      1
 0.15792824E+01 0.36528701E-03-0.50657672E-07-0.34884855E-10 0.88089699E-14    2
 0.99535752E+04-0.30240495E+01 0.58924019E+00 0.25012842E-02-0.34229498E-06    3
-0.18994346E-08 0.10190406E-11 0.10236923E+05 0.21937017E+01                   4
CH_Pt                  0C   1H   1PT  1     I    300.00   3000.00 1000.00      1
-0.48242472E-02 0.30446239E-02-0.16066099E-06-0.29041700E-09 0.57999924E-13    2
 0.22595219E+05 0.56677818E+01 0.84157485E+00 0.13095380E-02 0.28464575E-06    3
 0.63862904E-09-0.42766658E-12 0.22332801E+05 0.11452305E+01                   4
CH2_Pt                 0C   1H   2PT  1     I    300.00   3000.00 1000.00      1
 0.74076122E+00 0.48032533E-02-0.32825633E-06-0.47779786E-09 0.10073452E-12    2
 0.10443752E+05 0.40842086E+00-0.14876404E+00 0.51396289E-02 0.11211075E-05    3
-0.82755452E-09-0.44572345E-12 0.10878700E+05 0.57451882E+01                   4
CH3_Pt                 0C   1H   3PT  1     I    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
CO_Pt                  0C   1O   1PT  1     I    300.00   3000.00 1000.00      1
 0.47083778E+01 0.96037297E-03-0.11805279E-06-0.76883826E-10 0.18232000E-13    2
-0.32311723E+05-0.16719593E+02 0.48907466E+01 0.68134235E-04 0.19768814E-06    3
 0.12388669E-08-0.90339249E-12-0.32297836E+05-0.17453161E+02                   4
CO2_Pt            081292C   1O   2PT  1     I   300.00   3000.00  1000.00      1
 0.46900000E+00 0.62660000E-02 0.00000000E-00 0.00000000E-00 0.00000000E-00    2
-0.50458700E+05-0.45550000E+01 0.46900000E+00 0.62662000E-02 0.00000000E-00    3
 0.00000000E-00 0.00000000E-00-0.50458700E+05-0.45550000E+01                   4
H_Pt               92491H   1PT  1          I    300.00   3000.00 1000.00      1
 0.10696996E+01 0.15432230E-02-0.15500922E-06-0.16573165E-09 0.38359347E-13    2
-0.50546128E+04-0.71555238E+01-0.13029877E+01 0.54173199E-02 0.31277972E-06    3
-0.32328533E-08 0.11362820E-11-0.42277075E+04 0.58743238E+01                   4
H2O_Pt             92491O   1H   2PT  1     I    300.00   3000.00 1000.00      1
 0.25803051E+01 0.49570827E-02-0.46894056E-06-0.52633137E-09 0.11998322E-12    2
-0.38302234E+05-0.17406322E+02-0.27651553E+01 0.13315115E-01 0.10127695E-05    3
-0.71820083E-08 0.22813776E-11-0.36398055E+05 0.12098145E+02                   4
O_Pt               92491O   1PT  1          I    300.00   3000.00 1000.00      1
 0.19454180E+01 0.91761647E-03-0.11226719E-06-0.99099624E-10 0.24307699E-13    2
-0.14005187E+05-0.11531663E+02-0.94986904E+00 0.74042305E-02-0.10451424E-05    3
-0.61120420E-08 0.33787992E-11-0.13209912E+05 0.36137905E+01                   4
OH_Pt              92491O   1H   1PT  1     I    300.00   3000.00 1000.00      1
 0.18249973E+01 0.32501565E-02-0.31197541E-06-0.34603206E-09 0.79171472E-13    2
-0.26685492E+05-0.12280891E+02-0.20340881E+01 0.93662683E-02 0.66275214E-06    3
-0.52074887E-08 0.17088735E-11-0.25319949E+05 0.89863186E+01                   4
_Pt_                    PT  1               S    300.0    3000.0  1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
