!*******************************************************************************
! The following thermo data is from personal communication with 
! O. Deutschmann.  However, the reactions all have explicit reverse 
! reactions, so thermo data is not being used for reaction-rate calculations.
!*******************************************************************************

THERMO
   300.000  1000.000  5000.000
   
C3H6              120186C   3H   6          G  0300.00   5000.00  1000.00      1
 0.06732257E+02 0.14908336E-01-0.04949899E-04 0.07212022E-08-0.03766204E-12    2
-0.09235703E+04-0.13313348E+02 0.14933071E+01 0.02092517E+00 0.04486794E-04    3
-0.16689121E-07 0.07158146E-10 0.10748264E+04 0.16145340E+02                   4
H2                121286H   2               G   300.000  5000.000 1000.00      1
 2.99142300e+00 7.00064400e-04-5.63382900e-08-9.23157800e-12 1.58275200e-15    2
-8.35034000e+02-1.35511000e+00 3.29812400e+00 8.24944200e-04-8.14301500e-07    3
-9.47543400e-11 4.13487200e-13-1.01252100e+03-3.29409400e+00                   4
H2O                20387H   2O   1          G   300.000  5000.000 1000.00      1
 2.67214600e+00 3.05629300e-03-8.73026000e-07 1.20099600e-10-6.39161800e-15    2
-2.98992100e+04 6.86281700e+00 3.38684200e+00 3.47498200e-03-6.35469600e-06    3
 6.96858100e-09-2.50658800e-12-3.02081100e+04 2.59023300e+00                   4
CO                121286C   1O   1          G   300.000  5000.000 1000.00      1
 3.02507800e+00 1.44268900e-03-5.63082800e-07 1.01858100e-10-6.91095200e-15    2
-1.42683500e+04 6.10821800e+00 3.26245200e+00 1.51194100e-03-3.88175500e-06    3
 5.58194400e-09-2.47495100e-12-1.43105400e+04 4.84889700e+00                   4
CO2               121286C   1O   2          G   300.000  5000.000 1000.00      1
 4.45362300e+00 3.14016900e-03-1.27841100e-06 2.39399700e-10-1.66903300e-14    2
-4.89669600e+04-9.55395900e-01 2.27572500e+00 9.92207200e-03-1.04091100e-05    3
 6.86668700e-09-2.11728000e-12-4.83731400e+04 1.01884900e+01                   4
N2                121286N   2               G   300.000  5000.000 1000.00      1
 2.92664000e+00 1.48797700e-03-5.68476100e-07 1.00970400e-10-6.75335100e-15    2
-9.22797700e+02 5.98052800e+00 3.29867700e+00 1.40824000e-03-3.96322200e-06    3
 5.64151500e-09-2.44485500e-12-1.02090000e+03 3.95037200e+00                   4
NO                121286N   1O   1          G   300.000  5000.000 1000.00      1
 3.24543500e+00 1.26913800e-03-5.01589000e-07 9.16928300e-11-6.27541900e-15    2
 9.80084000e+03 6.41729400e+00 3.37654200e+00 1.25306300e-03-3.30275100e-06    3
 5.21781000e-09-2.44626300e-12 9.81796100e+03 5.82959000e+00                   4
O2                121386O   2               G   300.000  5000.000 1000.00      1
 3.69757800e+00 6.13519700e-04-1.25884200e-07 1.77528100e-11-1.13643500e-15    2
-1.23393000e+03 3.18916600e+00 3.21293600e+00 1.12748600e-03-5.75615000e-07    3
 1.31387700e-09-8.76855400e-13-1.00524900e+03 6.03473800e+00                   4

O(S)               92491O   1Pt  1          I    300.00   3000.00 1000.00      1
 0.19454180E+01 0.91761647E-03-0.11226719E-06-0.99099624E-10 0.24307699E-13    2
-0.14005187E+05-0.11531663E+02-0.94986904E+00 0.74042305E-02-0.10451424E-05    3
-0.61120420E-08 0.33787992E-11-0.13209912E+05 0.36137905E+01                   4
O2(S)              92491O   2Pt  1          I    300.00   3000.00 1000.00      1
 0.35989249E+01 0.20437732E-02-0.23878221E-06-0.22041054E-09 0.53299430E-13    2
-0.41095444E+04-0.21604582E+02-0.20174649E+01 0.14146218E-01-0.16376665E-05    3
-0.11264421E-07 0.60101386E-11-0.25084473E+04 0.79811935E+01                   4
H(S)               92491H   1Pt  1          I    300.00   3000.00 1000.00      1
 0.10696996E+01 0.15432230E-02-0.15500922E-06-0.16573165E-09 0.38359347E-13    2
-0.50546128E+04-0.71555238E+01-0.13029877E+01 0.54173199E-02 0.31277972E-06    3
-0.32328533E-08 0.11362820E-11-0.42277075E+04 0.58743238E+01                   4
H2(S)              92491H   2Pt  1          I    300.00   3000.00 1000.00      1
 0.15330955E+01 0.34586885E-02-0.32622225E-06-0.36824219E-09 0.83855205E-13    2
-0.36401533E+04-0.10822206E+02-0.21517782E+01 0.87039210E-02 0.11154106E-05    3
-0.42477102E-08 0.96133203E-12-0.22640681E+04 0.97397461E+01                   4
H2O(S)             92491O   1H   2Pt  1     I    300.00   3000.00 1000.00      1
 0.25803051E+01 0.49570827E-02-0.46894056E-06-0.52633137E-09 0.11998322E-12    2
-0.38302234E+05-0.17406322E+02-0.27651553E+01 0.13315115E-01 0.10127695E-05    3
-0.71820083E-08 0.22813776E-11-0.36398055E+05 0.12098145E+02                   4
OH(S)              92491O   1H   1Pt  1     I    300.00   3000.00 1000.00      1
 0.18249973E+01 0.32501565E-02-0.31197541E-06-0.34603206E-09 0.79171472E-13    2
-0.26685492E+05-0.12280891E+02-0.20340881E+01 0.93662683E-02 0.66275214E-06    3
-0.52074887E-08 0.17088735E-11-0.25319949E+05 0.89863186E+01                   4
Pt(S)                   Pt  1               S    300.0    3000.0  1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(S)                  0C   1O   1Pt  1     I    300.00   3000.00 1000.00      1
 0.47083778E+01 0.96037297E-03-0.11805279E-06-0.76883826E-10 0.18232000E-13    2
-0.32311723E+05-0.16719593E+02 0.48907466E+01 0.68134235E-04 0.19768814E-06    3
 0.12388669E-08-0.90339249E-12-0.32297836E+05-0.17453161E+02                   4
CO2(S)            081292C   1O   2Pt  1     I   300.00   3000.00  1000.00      1
 0.46900000E+00 0.62660000E-02 0.00000000E-00 0.00000000E-00 0.00000000E-00    2
-0.50458700E+05-0.45550000E+01 0.46900000E+00 0.62662000E-02 0.00000000E-00    3
 0.00000000E-00 0.00000000E-00-0.50458700E+05-0.45550000E+01                   4
C(S)                   0C   1Pt  1          I    300.00   3000.00 1000.00      1
 0.15792824E+01 0.36528701E-03-0.50657672E-07-0.34884855E-10 0.88089699E-14    2
 0.99535752E+04-0.30240495E+01 0.58924019E+00 0.25012842E-02-0.34229498E-06    3
-0.18994346E-08 0.10190406E-11 0.10236923E+05 0.21937017E+01                   4
CH(S)                  0C   1H   1Pt  1     I    300.00   3000.00 1000.00      1
-0.48242472E-02 0.30446239E-02-0.16066099E-06-0.29041700E-09 0.57999924E-13    2
 0.22595219E+05 0.56677818E+01 0.84157485E+00 0.13095380E-02 0.28464575E-06    3
 0.63862904E-09-0.42766658E-12 0.22332801E+05 0.11452305E+01                   4
CH2(S)                 0C   1H   2Pt  1     I    300.00   3000.00 1000.00      1
 0.74076122E+00 0.48032533E-02-0.32825633E-06-0.47779786E-09 0.10073452E-12    2
 0.10443752E+05 0.40842086E+00-0.14876404E+00 0.51396289E-02 0.11211075E-05    3
-0.82755452E-09-0.44572345E-12 0.10878700E+05 0.57451882E+01                   4
CH3(S)                 0C   1H   3Pt  1     I    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4
C3H6(S)                 C   3H   6Pt  2     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C3H5(S)                 C   3H   5Pt  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CC2H5(S)                C   3H   5Pt  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C2H3(S)                 C   2H   3Pt  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH3CO(S)                C   2H   3Pt  1O   1I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
NO(S)                   N   1O   1Pt  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
N(S)                    N   1Pt  1    0     I   300.0    3000.0   1000.        1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
NO2(S)                  N   1O   2Pt  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
Rh(S1)                  Rh  1               S   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
NO(S1)                  N   1O   1Rh  1     I   300.0    3000.0   1000.0       1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(S1)                 0C   1O   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
O(S1)              92491O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
N(S1)              92491N   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4

END
