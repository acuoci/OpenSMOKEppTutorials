!
! A. Stagni, C. Cavallotti, S. Arunthanayothin, Y. Song,
! O. Herbinet, F. Battin-Leclerc, T. Faravelli
! "An experimental, theoretical and kinetic-modeling study of the gas-phase oxidation of ammonia"
! Reaction Chemistry and Engineering (submitted) (2020).
!
! Submitted to Reaction Chemistry and Engineering (November 2019)
!
! Thermodynamic properties
! 
! CHEMKIN format
!
!VERSION:  17_03
!AUTHORS:  C1-C3   Burcat   
!NOTE:     SPECIES RE-ARRANGED AS THE SAME ORDER IN MECH
!
!VERSION:  17_05
!Following species are updated from ATcT's Database:
! H	H2	O	O2	HE
! OH	H2O	N2	HO2	HCO
! H2O2	AR	CO	CO2
 THERMO
  300.   1000.   4000.
!   ---------ARAMCO 2.0 -------------------
HE                ATcT3EHE  1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] He <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.49985609E+00 2.19365392E-07-1.07525085E-10 2.07198041E-14-1.39358612E-18    2
-7.45309155E+02 9.29535014E-01 2.49976293E+00 1.01013432E-06-8.24578465E-10    3
-6.85983306E-13 7.24751856E-16-7.45340917E+02 9.29800315E-01 0.00000000E+00    4
AR                ATcT3EAR  1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] Ar <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.49989176E+00 1.56134837E-07-7.76108557E-11 1.52928085E-14-1.05304493E-18    2
-7.45328403E+02 4.38029835E+00 2.49988611E+00 2.13037960E-07 8.97320772E-10    3
-2.31395752E-12 1.30201393E-15-7.45354481E+02 4.38024367E+00 0.00000000E+00    4
N2                ATcT3EN   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] N2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.93802970E+00 1.41838030E-03-5.03281045E-07 8.07555464E-11-4.76064275E-15    2
-9.17180990E+02 5.95521985E+00 3.53603521E+00-1.58270944E-04-4.26984251E-07    3
 2.37542590E-09-1.39708206E-12-1.04749645E+03 2.94603724E+00 0.00000000E+00    4
O2                ATcT3EO   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] O2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 3.65980488E+00 6.59877372E-04-1.44158172E-07 2.14656037E-11-1.36503784E-15    2
-1.21603048E+03 3.42074148E+00 3.78498258E+00-3.02002233E-03 9.92029171E-06    3
-9.77840434E-09 3.28877702E-12-1.06413589E+03 3.64780709E+00 0.00000000E+00    4
H2                ATcT3EH   2    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2 <g> ATcT ver. 1.122, DHf298 = 0.000 \B1 0.000 kJ/mol - fit MAR17
 2.90207649E+00 8.68992581E-04-1.65864430E-07 1.90851899E-11-9.31121789E-16    2
-7.97948726E+02-8.45591320E-01 2.37694204E+00 7.73916922E-03-1.88735073E-05    3
 1.95517114E-08-7.17095663E-12-9.21173081E+02 5.47184736E-01 0.00000000E+00    4
H2O               ATcT3EH   2O   1    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2O <g> ATcT ver. 1.122, DHf298 = -241.833 \B1 0.027 kJ/mol - fit MAR17
 2.73117512E+00 2.95136995E-03-8.35359785E-07 1.26088593E-10-8.40531676E-15    2
-2.99169082E+04 6.55183000E+00 4.20147551E+00-2.05583546E-03 6.56547207E-06    3
-5.52906960E-09 1.78282605E-12-3.02950066E+04-8.60610906E-01-2.90858262E+04    4
H2O2              ATcT3EH   2O   2    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H2O2 <g> ATcT ver. 1.122, DHf298 = -135.457 \B1 0.064 kJ/mol - fit MAR17
 4.54017480E+00 4.15970971E-03-1.30876777E-06 2.00823615E-10-1.15509243E-14    2
-1.79514029E+04 8.55881745E-01 4.23854160E+00-2.49610911E-04 1.59857901E-05    3
-2.06919945E-08 8.29766320E-12-1.76486003E+04 3.58850097E+00-1.62917334E+04    4
O                 ATcT3EO   1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] O <g> ATcT ver. 1.122, DHf298 = 249.229 \B1 0.002 kJ/mol - fit MAR17
 2.55160087E+00-3.83085457E-05 8.43197478E-10 4.01267136E-12-4.17476574E-16    2
 2.92287628E+04 4.87617014E+00 3.15906526E+00-3.21509999E-03 6.49255543E-06    3
-5.98755115E-09 2.06876117E-12 2.91298453E+04 2.09078344E+00 2.99753606E+04    4
H                 ATcT3EH   1    0    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] H <g> ATcT ver. 1.122, DHf298 = 217.998 \B1 0.000 kJ/mol - fit MAR17
 2.49985211E+00 2.34582548E-07-1.16171641E-10 2.25708298E-14-1.52992005E-18    2
 2.54738024E+04-4.45864645E-01 2.49975925E+00 6.73824499E-07 1.11807261E-09    3
-3.70192126E-12 2.14233822E-15 2.54737665E+04-4.45574009E-01 2.62191345E+04    4
OH                ATcT3EH   1O   1    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] OH <g> ATcT ver. 1.122, DHf298 = 37.490 \B1 0.027 kJ/mol - fit MAR17
 2.84581721E+00 1.09723818E-03-2.89121101E-07 4.09099910E-11-2.31382258E-15    2
 3.71706610E+03 5.80339915E+00 3.97585165E+00-2.28555291E-03 4.33442882E-06    3
-3.59926640E-09 1.26706930E-12 3.39341137E+03-3.55397262E-02 4.50901087E+03    4
HO2               ATcT3EH   1O   2    0    0G    200.00   6000.00 1000.00      1 ! [Ghobad] HO2 <g> ATcT ver. 1.122, DHf298 = 12.26 \B1 0.16 kJ/mol - fit MAR17 
 4.10564010E+00 2.04046836E-03-3.65877562E-07 1.85973044E-11 4.98818315E-16    2
 4.32898769E+01 3.30808126E+00 4.26251250E+00-4.45642032E-03 2.05164934E-05    3
-2.35794011E-08 9.05614257E-12 2.62442356E+02 3.88223684E+00 1.47417835E+03    4
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
!NOx MODULE (from Burcat http://garfield.chem.elte.hu/Burcat/THERM.DAT)
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NO                RUS 89N   1O   1    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.26071234E+00 1.19101135E-03-4.29122646E-07 6.94481463E-11-4.03295681E-15    2
 9.92143132E+03 6.36900518E+00 4.21859896E+00-4.63988124E-03 1.10443049E-05    3
-9.34055507E-09 2.80554874E-12 9.84509964E+03 2.28061001E+00 1.09770882E+04    4
N2O               L 7/88N   2O   1    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.48230729E+01 0.26270251E-02-0.95850872E-06 0.16000712E-09-0.97752302E-14    2
 0.80734047E+04-0.22017208E+01 0.22571502E+01 0.11304728E-01-0.13671319E-04    3
 0.96819803E-08-0.29307182E-11 0.87417746E+04 0.10757992E+02 0.98141682E+04    4
NO2               L 7/88N   1O   2    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.48847540E+01 0.21723955E-02-0.82806909E-06 0.15747510E-09-0.10510895E-13    2
 0.23164982E+04-0.11741695E+00 0.39440312E+01-0.15854290E-02 0.16657812E-04    3
-0.20475426E-07 0.78350564E-11 0.28966180E+04 0.63119919E+01 0.41124701E+04    4
HNO               ATcT/AH  1.N  1.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.16598124E+00 2.99958892E-03-3.94376786E-07-3.85344089E-11 7.07602668E-15    2
 1.17726311E+04 7.64511172E+00 4.53525574E+00-5.68543377E-03 1.85198540E-05    3
-1.71881225E-08 5.55818157E-12 1.16183003E+04 1.74315886E+00 1.28500657E+04    4
HNO2              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 4.66358504E+00 4.89854351E-03-1.79694193E-06 2.94420361E-10-1.78235577E-14    2
-7.25216334E+03-3.06053640E-02 4.03779347E+00-4.46123109E-03 3.19440815E-05    3
-3.79359490E-08 1.44570885E-11-6.53088236E+03 5.90620097E+00-5.31122753E+03    4
HONO              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 5.79144641E+00 3.64630732E-03-1.29112765E-06 2.06498233E-10-1.22138679E-14    2
-1.15974343E+04-4.07145349E+00 3.16416438E+00 8.50517773E-03 5.48561573E-07    3
-8.27656474E-09 4.39957151E-12-1.07744086E+04 1.00231941E+01-9.46242812E+03    4
HONO2             T 8/03H  1.N  1.O  3.   0.G   200.000  6000.000 1000.        1 ! HNO3 in Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 8.03098942E+00 4.46958589E-03-1.72459491E-06 2.91556153E-10-1.80102702E-14    2
-1.93138183E+04-1.62616537E+01 1.69329154E+00 1.90167702E-02-8.25176697E-06    3
-6.06113827E-09 4.65236978E-12-1.74198909E+04 1.71839838E+01-1.61524852E+04    4
N2H2      2/13/19       N   2H   2          G   300.000  5000.000 1380.000     1 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 4.14686796E+00 4.81612315E-03-1.62748817E-06 2.50556098E-10-1.44494188E-14    2
 2.33444055E+04 5.34122740E-01 2.55589425E+00 6.54339081E-03-8.81947855E-07    3
-1.15971304E-09 3.97442230E-13 2.41085081E+04 9.80504705E+00                   4
H2NN Isodiazene   T 9/11N  2.H  2.   0.   0.G   200.000  6000.000 1000.        1 ! Is 'N2H2 Isodiazene' in Burcat database
 3.05903670E+00 6.18382347E-03-2.22171165E-06 3.58539206E-10-2.14532905E-14    2
 3.48530149E+04 6.69893515E+00 4.53204001E+00-7.32418578E-03 3.00803713E-05    3
-3.04000551E-08 1.04700639E-11 3.49580003E+04 1.51074195E+00 3.61943157E+04    4
HNNO      5/30/18 THERM N  2.H  1.O  1    0.G   300.000  5000.000 1790.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 2.15594002E+06-4.13111192E+03 2.65627771E+00-6.70395293E-04 5.57827338E-08    2
-8.03468100E+08-1.18702032E+07-8.96779017E-01 3.69714359E-02-4.80099825E-05    3
 2.62274393E-08-5.11382966E-12 2.68675048E+04 2.64521806E+01                   4
NH2NO     5/30/18 THERM N  2.H  2.O  1    0.G   300.000  5000.000 1371.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 7.93898100E+00 5.21842622E-03-2.12493130E-06 3.53331059E-10-2.12447889E-14    2
 5.42322972E+03-1.84299492E+01 1.85914077E+00 1.68525394E-02-9.37240888E-06    3
 1.71380329E-09 4.84625807E-14 7.78108234E+03 1.51172833E+01                   4
HNOH trans & Equ  T11/11H  2.N  1.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.98321933E+00 4.88846374E-03-1.65086637E-06 2.55371446E-10-1.48308561E-14    2
 1.05780106E+04 3.62582838E+00 3.95608248E+00-3.02611020E-03 2.56874396E-05    3
-3.15645120E-08 1.24084574E-11 1.09199790E+04 5.55950983E+00 1.21354115E+04    4
NH2OH             ATcT/AN  1.H  3.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.88112502E+00 8.15708448E-03-2.82615576E-06 4.37930933E-10-2.52724604E-14    2
-6.86018419E+03 3.79156136E+00 3.21016092E+00 6.19671676E-03 1.10594948E-05    3
-1.96668262E-08 8.82516590E-12-6.58148481E+03 7.93293571E+00-5.28593988E+03    4
NH3               ATcT3EH   3N   1    0    0G    200.00   4000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 2.36074311E+00 6.31850146E-03-2.28966806E-06 4.11767411E-10-2.90836787E-14    2
-6.41596473E+03 8.02154329E+00 4.14027871E+00-3.58489142E-03 1.89475904E-05    3
-1.98833970E-08 7.15267961E-12-6.68545158E+03-1.66754883E-02-5.47888720E+03    4
N2H4 HYDRAZINE    L 5/90N   2H   4    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 4.93957357E+00 8.75017187E-03-2.99399058E-06 4.67278418E-10-2.73068599E-14    2
 9.28265548E+03-2.69439772E+00 3.83472149E+00-6.49129555E-04 3.76848463E-05    3
-5.00709182E-08 2.03362064E-11 1.00893925E+04 5.75272030E+00 1.14474575E+04    4
N                 L 6/88N   1    0    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.24159429E+01 0.17489065E-03-0.11902369E-06 0.30226244E-10-0.20360983E-14    2
 0.56133775E+05 0.46496095E+01 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.56104638E+05 0.41939088E+01 0.56850013E+05    4
NO3               ATcT/AN  1.O  3.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 7.48347702E+00 2.57772064E-03-1.00945831E-06 1.72314063E-10-1.07154008E-14    2
 6.12990474E+03-1.41618136E+01 2.17359330E+00 1.04902685E-02 1.10472669E-05    3
-2.81561867E-08 1.36583960E-11 7.81290905E+03 1.46022090E+01 8.97563416E+03    4
NH                ATcT/AN  1.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 2.78372644E+00 1.32985888E-03-4.24785573E-07 7.83494442E-11-5.50451310E-15    2
 4.23461945E+04 5.74084863E+00 3.49295037E+00 3.11795720E-04-1.48906628E-06    3
 2.48167402E-09-1.03570916E-12 4.21059722E+04 1.84834973E+00 4.31525130E+04    4
NNH               T 8/11N  2.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! N2H in Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.42744423E+00 3.23295234E-03-1.17296299E-06 1.90508356E-10-1.14491506E-14    2
 2.87676026E+04 6.39209233E+00 4.25474632E+00-3.45098298E-03 1.37788699E-05    3
-1.33263744E-08 4.41023397E-12 2.87932080E+04 3.28551762E+00 3.00058572E+04    4
NH2  AMIDOGEN RAD IU3/03N  1.H  2.   0.   0.G   200.000  3000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 2.59263049E+00 3.47683597E-03-1.08271624E-06 1.49342558E-10-5.75241187E-15    2
 2.15737320E+04 7.90565351E+00 4.19198016E+00-2.04602827E-03 6.67756134E-06    3
-5.24907235E-09 1.55589948E-12 2.11863286E+04-9.04785244E-02 2.23945849E+04    4
H2NO  RADICAL     T09/09N  1.H  2.O  1.   0.G   200.000  6000.000 1000.        1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 3.75555914E+00 5.16219354E-03-1.76387387E-06 2.75052692E-10-1.60643143E-14    2
 6.51826177E+03 4.30933053E+00 3.93201139E+00-1.64028165E-04 1.39161409E-05    3
-1.62747853E-08 6.00352834E-12 6.71178975E+03 4.58837038E+00 7.97044877E+03    4
N2H3   Rad.       T 7/11N  2.H  3.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 4.04483566E+00 7.31130186E-03-2.47625799E-06 3.83733021E-10-2.23107573E-14    2
 2.53241420E+04 2.88423392E+00 3.42125505E+00 1.34901590E-03 2.23459071E-05    3
-2.99727732E-08 1.20978970E-11 2.58198956E+04 7.83176309E+00 2.70438066E+04    4
END
