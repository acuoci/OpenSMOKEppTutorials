!***********************************************************************
!****     CO/O2 OVER RH - SURFASE MECHANISM                            *
!****     thermodynamically constant (273 - 1273K)                     *
!****                                                                  *
!****     References:                                                  *
!****     H. Karadeniz, C. Karakaya, S. Tischer, O. Deutschmann,       *
!****     Chemical Engineering Science, Submitted (2013).              *
!****     www.detchem.com/mechanisms                                   * 
!****     KIT (Karlsruhe Institute of Technology)                      *
!****     Contact: mail@detchem.com (O. Deutschmann)                   * 
!****     www.detchem.com/mechanisms                                   * 
!****                                                                  *
!****                                                                  *
!****     Kinetic data:                                                *
!****      k = A * T**b * exp (-Ea/RT)         A          b       Ea   *
!****                                       (cm,mol,s)    -     kJ/mol *
!****                                                                  *
!****     STICK: A in next reaction is initial sticking coefficient    *
!****                                                                  *
!****                                                                  *
!****     (CHEMKIN format)                                             *
!****                                                                  * 
!***********************************************************************     

THERMO
   300.000  1000.000  3000.000

AR            (adjust)  AR  1    0    0    0G   300.00   5000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
N2                      N   2    0    0    0G   300.00   5000.00  1000.00      1
 2.85328990E+00 1.60221280E-03-6.29368930E-07 1.14410220E-10-7.80574650E-15    2
-8.90080930E+02 6.39648970E+00 3.70441770E+00-1.42187530E-03 2.86703920E-06    3
-1.20288850E-09-1.39546770E-14-1.06407950E+03 2.23362850E+00                   4
O(s)                    O   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
O2(s)                   O   2Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H(s)                    H   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2(s)                   H   2Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O(s)                  O   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
OH(s)                   O   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
Rh(s)                   Rh  1               S    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO(s)                   C   1O   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CO2(s)                  C   1O   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
C(s)                    C   1Rh  1          I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH(s)                   C   1H   1Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH2(s)                  C   1H   2Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH3(s)                  C   1H   3Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH4(s)                  C   1H   4Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
HCO(s)                  C   1H   1Rh  1O   1I    300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
CH4           (adjust)  C   1H   4    0    0     300.00   5000.00 1000.00      1
 1.68347883E+00 1.02372356E-02-3.87512864E-06 6.78558487E-10-4.50342312E-14    2
-1.00807871E+04 9.62339497E+00 7.78741479E-01 1.74766835E-02-2.78340904E-05    3
 3.04970804E-08-1.22393068E-11-9.82522852E+03 1.37221947E+01                   4
O2            (adjust)  O   2    0    0    0     300.00   5000.00 1000.00      1
 3.61221390E+00 7.48531660E-04-1.98206470E-07 3.37490080E-11-2.39073740E-15    2
-1.19781510E+03 3.67033070E+00 3.78371350E+00-3.02336340E-03 9.94927510E-06    3
-9.81891010E-09 3.30318250E-12-1.06381070E+03 3.64163450E+00                   4
CO            (adjust)  C   1O   1    0    0     300.00   5000.00 1000.00      1
 3.02507806E+00 1.44268852E-03-5.63082779E-07 1.01858133E-10-6.91095156E-15    2
-1.42683496E+04 6.10821772E+00 3.26245165E+00 1.51194085E-03-3.88175522E-06    3
 5.58194424E-09-2.47495123E-12-1.43105391E+04 4.84889698E+00                   4
CO2           (adjust)  C   1O   2    0    0     300.00   5000.00 1000.00      1
 4.45362282E+00 3.14016873E-03-1.27841054E-06 2.39399667E-10-1.66903319E-14    2
-4.89669609E+04-9.55395877E-01 2.27572465E+00 9.92207229E-03-1.04091132E-05    3
 6.86668678E-09-2.11728009E-12-4.83731406E+04 1.01884880E+01                   4
H2            (adjust)  H   2    0    0    0     300.00   5000.00 1000.00      1
 3.06670950E+00 5.74737550E-04 1.39383190E-08-2.54835180E-11 2.90985740E-15    2
-8.65474120E+02-1.77984240E+00 3.35535140E+00 5.01361440E-04-2.30069080E-07    3
-4.79053240E-10 4.85225850E-13-1.01916260E+03-3.54772280E+00                   4
H2O           (adjust)  H   2O   1    0    0     300.00   5000.00 1000.00      1
 2.61104720E+00 3.15631300E-03-9.29854380E-07 1.33315380E-10-7.46893510E-15    2
-2.98681670E+04 7.20912680E+00 4.16772340E+00-1.81149700E-03 5.94712880E-06    3
-4.86920210E-09 1.52919910E-12-3.02899690E+04-7.31354740E-01                   4
AR            (adjust)  AR  1    0    0    0     300.00   5000.00 1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375020E+02 4.36600060E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45374980E+02 4.36600060E+00                   4
NI(*)         (adjust)  NI  1    0    0    0     300.00   3000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
H2O(*)        (adjust)  H   2O   1NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-3.28621348E+04 1.57219174E+01 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-3.28621348E+04 1.57219174E+01                   4
H(*)          (adjust)  H   1NI  1    0    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-3.82656399E+03 4.89898398E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-3.82656399E+03 4.89898398E+00                   4
COOH(*)       (adjust)  C   1H   1O   2NI  1     300.00   5000.00 1000.00      1
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00                   4
OH(*)         (adjust)  H   1O   1NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-2.31833113E+04 1.28038592E+01 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-2.31833113E+04 1.28038592E+01                   4
CO(*)         (adjust)  C   1O   1NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-2.37539453E+04 1.96355620E+01 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-2.37539453E+04 1.96355620E+01                   4
C(*)          (adjust)  C   1NI  1    0    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-9.60170600E+02-9.94267012E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-9.60170600E+02-9.94267012E+00                   4
CH3(*)        (adjust)  C   1H   3NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-3.58843376E+03 3.36230167E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-3.58843376E+03 3.36230167E+00                   4
CH2(*)        (adjust)  C   1H   2NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 5.94161025E+03 2.12413716E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 5.94161025E+03 2.12413716E+00                   4
CH(*)         (adjust)  C   1H   1NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 1.22543876E+04-2.56790500E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 1.22543876E+04-2.56790500E+00                   4
CH4(*)        (adjust)  C   1H   4NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.27928907E+03 8.44319611E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.27928907E+03 8.44319611E+00                   4
O(*)          (adjust)  O   1NI  1    0    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-2.66580549E+04 4.68860658E+00 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-2.66580549E+04 4.68860658E+00                   4
CO2(*)        (adjust)  C   1O   2NI  1    0     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-4.59500678E+04 2.14541635E+01 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-4.59500678E+04 2.14541635E+01                   4
HCO(*)        (adjust)  C   1H   1O   1NI  1     293.00   5000.00 5000.00      1
 1.00000000E-99 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-1.21882034E+04 1.49580180E+01 1.00000000E-99 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-1.21882034E+04 1.49580180E+01                   4
C3H8(s)       (adjust)  C   3H   8Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
C2H3(s)       (adjust)  C   2H   3Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
C3H7(s)       (adjust)  C   3H   7Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
C3H6(s)       (adjust)  C   3H   6Rh  1     I    300.00   3000.00 1000.00      1
 0.00000000E-00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-0.00000000E+00-0.00000000E+00 0.00000000E-00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-0.00000000E+00-0.00000000E+00                   4
C3H8              120186C   3H   8          G  0300.00   5000.00  1000.00      1
 0.07525217E+02 0.01889034E+00-0.06283924E-04 0.09179373E-08-0.04812410E-12    2
-0.16464548E+05-0.01784390E+03 0.08969208E+01 0.02668986E+00 0.05431425E-04    3
-0.02126000E-06 0.09243330E-10-0.13954918E+05 0.01935533E+03                   4
COOH(s)                 C   1H   1O   2Rh  1I    300.00   3000.00 1000.00      1
 0.30016165E+01 0.54084505E-02-0.40538058E-06-0.53422466E-09 0.11451887E-12    2
-0.32752722E+04-0.10965984E+02 0.12919217E+01 0.72675603E-02 0.98179476E-06    3
-0.20471294E-08 0.90832717E-13-0.25745610E+04-0.11983037E+01                   4

END
